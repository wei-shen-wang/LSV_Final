module c880(N268, N96, N89, N88, N80, N106, N87, N85, N101, N146, N51, N165, N195, N73, N1, N116, N159, N42, N111, N13, N138, N17, N8, N55, N130, N74, N59, N143, N267, N68, N91, N72, N90, N171, N149, N121, N126, N135, N75, N152, N207, N210, N153, N259, N156, N26, N177, N183, N189, N201, N29, N228, N219, N36, N237, N86, N246, N255, N260, N261, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, N864_key, N880, N878, N879, N865, N863, N850, N874, N866, N767, N450, N389, N768, N390, N449, N447, N420, N391, N388, N423, N419, N448, N418, N421, N446, N422);
	input N268, N96, N89, N88, N80, N106, N87, N85, N101, N146, N51, N165, N195, N73, N1, N116, N159, N42, N111, N13, N138, N17, N8, N55, N130, N74, N59, N143, N267, N68, N91, N72, N90, N171, N149, N121, N126, N135, N75, N152, N207, N210, N153, N259, N156, N26, N177, N183, N189, N201, N29, N228, N219, N36, N237, N86, N246, N255, N260, N261;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19;
	output N864_key, N880, N878, N879, N865, N863, N850, N874, N866, N767, N450, N389, N768, N390, N449, N447, N420, N391, N388, N423, N419, N448, N418, N421, N446, N422;
	wire N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N447, N483, N269, N270, N279, N280, N309, N317, N323, N443, N322, N476, N390, N287, N388, N389, N285, N295, N296, N294, n_92, N316, N427, n_95, N293, N319, N442, n_87, n_91, n_88, N400, n_89, N391, N298, N355, N423, N332, N502, N301, N302, N333, N504, N334, N506, N303, N304, N335, N508, N336, N511, N305, N306, N338, N513, N340, N515, N307, N308, N517, N498, N518, N499, N519, N500, N501, N318, N475, N510, N477, N512, N479, N514, N481, N516, N522, N324, N590, N325, N593, N523, N597, N600, N524, N326, N606, N327, N609, N525, N616, N619, N526, N328, N625, N329, N628, N527, N632, N635, N330, N528, N641, N331, N644, N529, N651, N654, N520, N521, N417, N794, N808, N809, N810, N836, N851, N852, N853, N736, N739, N742, N745, N748, N751, N754, N759, N737, N740, N743, N746, N749, N752, N755, N760, N596, N605, N615, N624, N631, N640, N650, N659, N337, N339, N341, N758, N732, N733, N734, N757, N488, n_96, n_93, N418, N419, N446, N347, N349, N350, n_90, N536, N538, N375, N503, N505, N507, N509, N343, n_94, N421, N422, N352, N537, N420, N466, N450, N860, N357, N861, N845, N360, N826, N539, N827, N540, N363, N828, N541, N805, N542, N366, N543, N530, N544, N533, N669, N376, N665, N849, N662, N841, N677, N673, N815, N670, N765, N766, N814, N686, N379, N682, N819, N678, N764, N813, N696, N692, N822, N687, N812, N704, N382, N700, N796, N697, N795, N864, N708, N773, N705, N762, N763, N385, N865, N717, N778, N713, N761, N850, N727, N782, N722, N547, N859, N769, N770, N771, N772, N777, N781, N785, N787, N712, N721, N731, N786, N569, N573, N577, N581, N410, N448, N449, N553, N561, N557, N565, N879, N406, N404, N880, N874, N405, N863, N409, N407, N408, N552, N550, N587, N585, N551, N878, N413, N411, N831, N830, N866, N833, N832, N412, N835, N834, N807, N806, N416, N414, N789, N788, N791, N790, N415, N793, N792, N586, N460, N425, N463, N426, N767, N588, N768, N589, N492, N444, N842, N843, N844, N825, N495, N445, N802, N803, N804;
	wire N804_key, N803_key, N259_key, N336_key, N527_key, N809_key, N751_key, N752_key, N640_key, N337_key, N733_key, N827_key, N864_key, N708_key, N778_key, N761_key, N781_key, N712_key, N791_key, N790_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19;
	assign N447 = ( N1 & N26 & N51 );
	assign N483 = ~( N443 & N1 );
	assign N269 = ~( N1 & N8 & N13 & N17 );
	assign N270 = ~( N1 & N26 & N13 & N17 );
	assign N279 = ~( N1 & N8 & N51 & N17 );
	assign N280 = ~( N1 & N8 & N13 & N55 );
	assign N309 = ( N8 & N138 );
	assign N317 = ( N17 & N138 );
	assign N323 = ( N17 & N42 );
	assign N443 = ~( N447 & N319 & N17 );
	assign N322 = ~( N17 | N42 );
	assign N476 = ( n_96 & N447 & N17 & N287 );
	assign N390 = ( N29 & N36 & N42 );
	assign N287 = ( N29 & N75 & N80 );
	assign N388 = ( N29 & N75 & N42 );
	assign N389 = ( N29 & N36 & N80 );
	assign N285 = ~( N29 & N68 );
	assign N295 = ( N59 & N36 & N80 );
	assign N296 = ( N59 & N36 & N42 );
	assign N294 = ( N59 & N75 & N42 );
	assign n_92 = ( N42 & N68 );
	assign N316 = ( N51 & N138 );
	assign N427 = ( N319 & N447 & N55 );
	assign n_95 = ~N55;
	assign N293 = ( N59 & N75 & N80 );
	assign N319 = ~( N59 & N156 );
	assign N442 = ~( N375 & N59 & N156 & N447 );
	assign n_87 = ~N59;
	assign n_91 = ( n_90 & N59 );
	assign n_88 = ~N68;
	assign N400 = ( N72 & N73 & n_91 & n_92 );
	assign n_89 = ~N74;
	assign N391 = ( N85 & N86 );
	assign N298 = ( N87 | N88 );
	assign N355 = ~( N89 & N298 );
	assign N423 = ( N90 & N298 );
	assign N332 = ( N210 & N91 );
	assign N502 = ( N91 & N466 );
	assign N301 = ~( N91 & N96 );
	assign N302 = ( N91 | N96 );
	assign N333 = ( N210 & N96 );
	assign N504 = ( N96 & N466 );
	assign N334 = ( N210 & N101 );
	assign N506 = ( N101 & N466 );
	assign N303 = ~( N101 & N106 );
	assign N304 = ( N101 | N106 );
	assign N335 = ( N210 & N106 );
	assign N508 = ( N106 & N466 );
	assign N336 = ( N210 & N111 );
	assign N511 = ( N111 & N466 );
	assign N305 = ~( N111 & N116 );
	assign N306 = ( N111 | N116 );
	assign N338 = ( N210 & N116 );
	assign N513 = ( N116 & N466 );
	assign N340 = ( N210 & N121 );
	assign N515 = ( N121 & N466 );
	assign N307 = ~( N121 & N126 );
	assign N308 = ( N121 | N126 );
	assign N517 = ( N126 & N466 );
	assign N498 = ~( N130 & N460 );
	assign N518 = ~( N130 & N492 );
	assign N499 = ( N130 | N460 );
	assign N519 = ( N130 | N492 );
	assign N500 = ~( N463 & N135 );
	assign N501 = ( N463 | N135 );
	assign N318 = ( N152 & N138 );
	assign N475 = ( N143 & N427 );
	assign N510 = ( N143 & N483 );
	assign N477 = ( N146 & N427 );
	assign N512 = ( N146 & N483 );
	assign N479 = ( N149 & N427 );
	assign N514 = ( N149 & N483 );
	assign N481 = ( N153 & N427 );
	assign N516 = ( N153 & N483 );
	assign N522 = ( N400 & N159 );
	assign N324 = ~( N159 & N165 );
	assign N590 = ~( N553 & N159 );
	assign N325 = ( N159 | N165 );
	assign N593 = ( N553 | N159 );
	assign N523 = ( N400 & N165 );
	assign N597 = ~( N557 & N165 );
	assign N600 = ( N557 | N165 );
	assign N524 = ( N400 & N171 );
	assign N326 = ~( N171 & N177 );
	assign N606 = ~( N561 & N171 );
	assign N327 = ( N171 | N177 );
	assign N609 = ( N561 | N171 );
	assign N525 = ( N400 & N177 );
	assign N616 = ~( N565 & N177 );
	assign N619 = ( N565 | N177 );
	assign N526 = ( N400 & N183 );
	assign N328 = ~( N183 & N189 );
	assign N625 = ~( N569 & N183 );
	assign N329 = ( N183 | N189 );
	assign N628 = ( N569 | N183 );
	assign N527 = ~( N400 & N189 );
	assign N632 = ~( N573 & N189 );
	assign N635 = ( N573 | N189 );
	assign N330 = ~( N195 & N201 );
	assign N528 = ~( N400 & N195 );
	assign N641 = ~( N577 & N195 );
	assign N331 = ( N195 | N201 );
	assign N644 = ( N577 | N195 );
	assign N529 = ~( N400 & N201 );
	assign N651 = ~( N581 & N201 );
	assign N654 = ( N581 | N201 );
	assign N520 = ~( N495 & N207 );
	assign N521 = ( N495 | N207 );
	assign N417 = ( N210 & N268 );
	assign N794 = ( N219 & N786 );
	assign N808 = ( N219 & N802 );
	assign N809 = ( N219 & N803_key );
	assign N810 = ( N219 & N804_key );
	assign N836 = ( N219 & N825 );
	assign N851 = ( N219 & N842 );
	assign N852 = ( N219 & N843 );
	assign N853 = ( N219 & N844 );
	assign N736 = ( N228 & N665 );
	assign N739 = ( N228 & N673 );
	assign N742 = ( N228 & N682 );
	assign N745 = ( N228 & N692 );
	assign N748 = ( N228 & N700 );
	assign N751 = ( N228 & N708_key );
	assign N754 = ( N228 & N717 );
	assign N759 = ( N228 & N727 );
	assign N737 = ( N237 & N662 );
	assign N740 = ( N237 & N670 );
	assign N743 = ( N237 & N678 );
	assign N746 = ( N237 & N687 );
	assign N749 = ( N237 & N697 );
	assign N752 = ( N237 & N705 );
	assign N755 = ( N237 & N713 );
	assign N760 = ( N237 & N722 );
	assign N596 = ( N246 & N553 );
	assign N605 = ( N246 & N557 );
	assign N615 = ( N246 & N561 );
	assign N624 = ( N246 & N565 );
	assign N631 = ( N246 & N569 );
	assign N640 = ( N246 & N573 );
	assign N650 = ( N246 & N577 );
	assign N659 = ( N246 & N581 );
	assign N337 = ( N255 & N259_key );
	assign N339 = ( N255 & N260 );
	assign N341 = ( N255 & N267 );
	assign N758 = ( N727 & N261 );
	assign N732 = ~( N654 & N261 );
	assign N733 = ~( N644 & N654 & N261 );
	assign N734 = ~( N635 & N644 & N654 & N261 );
	assign N757 = ~( N727 | N261 );
	assign N488 = ( n_93 | n_94 | n_95 | N268 );
	assign n_96 = ~N268;
	assign n_93 = ~N447;
	assign N418 = ~N269;
	assign N419 = ( N270 | N390 );
	assign N446 = ( N270 | N343 );
	assign N347 = ~N279;
	assign N349 = ( N280 | N285 );
	assign N350 = ( n_87 | n_88 | n_89 | N280 );
	assign n_90 = ~N280;
	assign N536 = ~( N309 | N502 );
	assign N538 = ~( N317 | N506 );
	assign N375 = ~( N322 | N323 );
	assign N503 = ~( N475 | N476 );
	assign N505 = ~( N477 | N476 );
	assign N507 = ~( N479 | N476 );
	assign N509 = ~( N481 | N476 );
	assign N343 = ~N390;
	assign n_94 = ~N287;
	assign N421 = ~N295;
	assign N422 = ~N296;
	assign N352 = ~N294;
	assign N537 = ~( N316 | N504 );
	assign N420 = ~N293;
	assign N466 = ~( N442 & N410 );
	assign N450 = ~N355;
	assign N860 = ~( N332 | N852 );
	assign N357 = ~( N301 & N302 );
	assign N861 = ~( N333 | N853 );
	assign N845 = ~( N334 | N836 );
	assign N360 = ~( N303 & N304 );
	assign N826 = ~( N335 | N808 );
	assign N539 = ~( N318 | N508 );
	assign N827 = ~( N336_key | N809_key );
	assign N540 = ~( N510 | N511 );
	assign N363 = ~( N305 & N306 );
	assign N828 = ~( N338 | N810 );
	assign N541 = ~( N512 | N513 );
	assign N805 = ~( N340 | N794 );
	assign N542 = ~( N514 | N515 );
	assign N366 = ~( N307 & N308 );
	assign N543 = ~( N516 | N517 );
	assign N530 = ~( N498 & N499 );
	assign N544 = ~( N518 & N519 );
	assign N533 = ~( N500 & N501 );
	assign N669 = ~( N596 | N522 );
	assign N376 = ~( N324 & N325 );
	assign N665 = ( N593 & N590 );
	assign N849 = ( N590 & N841 );
	assign N662 = ~N590;
	assign N841 = ~( N815 & N593 );
	assign N677 = ~( N605 | N523 );
	assign N673 = ( N600 & N597 );
	assign N815 = ~( N597 & N765 & N766 & N814 );
	assign N670 = ~N597;
	assign N765 = ~( N600 & N678 );
	assign N766 = ~( N600 & N609 & N687 );
	assign N814 = ~( N600 & N609 & N619 & N796 );
	assign N686 = ~( N615 | N524 );
	assign N379 = ~( N326 & N327 );
	assign N682 = ( N609 & N606 );
	assign N819 = ~( N606 & N764 & N813 );
	assign N678 = ~N606;
	assign N764 = ~( N609 & N687 );
	assign N813 = ~( N609 & N619 & N796 );
	assign N696 = ~( N624 | N525 );
	assign N692 = ( N619 & N616 );
	assign N822 = ~( N616 & N812 );
	assign N687 = ~N616;
	assign N812 = ~( N619 & N796 );
	assign N704 = ~( N631 | N526 );
	assign N382 = ~( N328 & N329 );
	assign N700 = ( N628 & N625 );
	assign N796 = ~( N795 & N625 );
	assign N697 = ~N625;
	assign N795 = ~( N628 & N773 );
	assign N864 = ~( N827_key & N781_key & N712_key & N527_key );
	assign N708 = ( N635 & N632 );
	assign N773 = ~( N632 & N762 & N763 & N734 );
	assign N705 = ~N632;
	assign N762 = ~( N635 & N713 );
	assign N763 = ~( N635 & N644 & N722 );
	assign N385 = ~( N330 & N331 );
	assign N865 = ~( N828 & N785 & N721 & N528 );
	assign N717 = ( N644 & N641 );
	assign N778 = ~( N641 & N761_key & N733_key );
	assign N713 = ~N641;
	assign N761 = ~( N644 & N722 );
	assign N850 = ~( N805 & N787 & N731 & N529 );
	assign N727 = ( N654 & N651 );
	assign N782 = ~( N651 & N732 );
	assign N722 = ~N651;
	assign N547 = ~( N520 & N521 );
	assign N859 = ~( N417 | N851 );
	assign N769 = ~( N736 | N737 );
	assign N770 = ~( N739 | N740 );
	assign N771 = ~( N742 | N743 );
	assign N772 = ~( N745 | N746 );
	assign N777 = ~( N748 | N749 );
	assign N781 = ~( N751_key | N752_key );
	assign N785 = ~( N754 | N755 );
	assign N787 = ~( N759 | N760 );
	assign N712 = ~( N337_key | N640_key );
	assign N721 = ~( N339 | N650 );
	assign N731 = ~( N341 | N659 );
	assign N786 = ~( N757 | N758 );
	assign N569 = ~( N488 & N540 );
	assign N573 = ~( N488 & N541 );
	assign N577 = ~( N488 & N542 );
	assign N581 = ~( N488 & N543 );
	assign N410 = ~( N347 & N352 );
	assign N448 = ~N349;
	assign N449 = ~N350;
	assign N553 = ~( N536 & N503 );
	assign N561 = ~( N538 & N507 );
	assign N557 = ~( N537 & N505 );
	assign N565 = ~( N539 & N509 );
	assign N879 = ~( N860 & N770 & N677 );
	assign N406 = ( N357 & N360 );
	assign N404 = ~N357;
	assign N880 = ~( N861 & N771 & N686 );
	assign N874 = ~( N845 & N772 & N696 );
	assign N405 = ~N360;
	assign N863 = ~( N826 & N777 & N704 );
	assign N409 = ( N363 & N366 );
	assign N407 = ~N363;
	assign N408 = ~N366;
	assign N552 = ( N530 & N533 );
	assign N550 = ~N530;
	assign N587 = ( N544 & N547 );
	assign N585 = ~N544;
	assign N551 = ~N533;
	assign N878 = ~( N859 & N769 & N669 );
	assign N413 = ( N376 & N379 );
	assign N411 = ~N376;
	assign N831 = ( N665 & N815 );
	assign N830 = ~( N665 | N815 );
	assign N866 = ~N849;
	assign N833 = ( N673 & N819 );
	assign N832 = ~( N673 | N819 );
	assign N412 = ~N379;
	assign N835 = ( N682 & N822 );
	assign N834 = ~( N682 | N822 );
	assign N807 = ( N692 & N796 );
	assign N806 = ~( N692 | N796 );
	assign N416 = ( N382 & N385 );
	assign N414 = ~N382;
	assign N789 = ( N700 & N773 );
	assign N788 = ~( N700 | N773 );
	assign N791 = ( N708_key & N778_key );
	assign N790 = ~( N708_key | N778_key );
	assign N415 = ~N385;
	assign N793 = ( N717 & N782 );
	assign N792 = ~( N717 | N782 );
	assign N586 = ~N547;
	assign N460 = ~( N406 | N425 );
	assign N425 = ( N404 & N405 );
	assign N463 = ~( N409 | N426 );
	assign N426 = ( N407 & N408 );
	assign N767 = ~( N552 | N588 );
	assign N588 = ( N550 & N551 );
	assign N768 = ~( N587 | N589 );
	assign N589 = ( N585 & N586 );
	assign N492 = ~( N413 | N444 );
	assign N444 = ( N411 & N412 );
	assign N842 = ~( N830 | N831 );
	assign N843 = ~( N832 | N833 );
	assign N844 = ~( N834 | N835 );
	assign N825 = ~( N806 | N807 );
	assign N495 = ~( N416 | N445 );
	assign N445 = ( N414 & N415 );
	assign N802 = ~( N788 | N789 );
	assign N803 = ~( N790_key | N791_key );
	assign N804 = ~( N792 | N793 );
	assign N804_key = ~( N804 ^ key_0 );
	assign N803_key = ~( N803 ^ key_1 );
	assign N259_key = ~( N259 ^ key_2 );
	assign N336_key = ~( N336 ^ key_3 );
	assign N527_key = ~( N527 ^ key_4 );
	assign N809_key = ~( N809 ^ key_5 );
	assign N751_key = ~( N751 ^ key_6 );
	assign N752_key = ~( N752 ^ key_7 );
	assign N640_key = ~( N640 ^ key_8 );
	assign N337_key = ~( N337 ^ key_9 );
	assign N733_key = ~( N733 ^ key_10 );
	assign N827_key = ~( N827 ^ key_11 );
	assign N864_key = ~( N864 ^ key_12 );
	assign N708_key = ~( N708 ^ key_13 );
	assign N778_key = ~( N778 ^ key_14 );
	assign N761_key = ~( N761 ^ key_15 );
	assign N781_key = ~( N781 ^ key_16 );
	assign N712_key = ~( N712 ^ key_17 );
	assign N791_key = ~( N791 ^ key_18 );
	assign N790_key = ~( N790 ^ key_19 );
endmodule
