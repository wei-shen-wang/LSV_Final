module c1908(N104, N91, N37, N31, N46, N79, N25, N10, N19, N13, N22, N43, N4, N49, N56, N99, N1, N63, N40, N34, N53, N16, N72, N60, N66, N82, N69, N94, N85, N7, N76, N28, N88, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, N2892, N2891, N2890, N2888, N2887, N2886, N2787, N2889, N2785, N2753, N2782, N2755, N2811, N2762, N2754, N2756, N2767, N2768, N2779, N2783, N2780, N2899, N2781, N2786, N2784);
	input N104, N91, N37, N31, N46, N79, N25, N10, N19, N13, N22, N43, N4, N49, N56, N99, N1, N63, N40, N34, N53, N16, N72, N60, N66, N82, N69, N94, N85, N7, N76, N28, N88;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25;
	output N2892, N2891, N2890, N2888, N2887, N2886, N2787, N2889, N2785, N2753, N2782, N2755, N2811, N2762, N2754, N2756, N2767, N2768, N2779, N2783, N2780, N2899, N2781, N2786, N2784;
	wire N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88, N91, N94, N99, N104, N1160, N1443, N2720, N190, N1309, N1387, N2721, N194, N1206, N1397, N2722, N197, N1054, N1226, N1345, N2723, N201, N1119, N1447, N2757, N206, N1128, N1311, N2758, N209, N1132, N1210, N2759, N212, N1055, N1120, N1129, N2760, N216, N1063, N1678, N2761, N220, N1130, N1133, N1453, N2734, N225, N1389, N1457, N2763, N229, N1315, N1399, N2764, N232, N1067, N1221, N2765, N235, N1064, N1317, N2766, N239, N1122, N1131, N1313, N2743, N243, N1214, N1462, N2744, N247, N592, N907, N2812, N724, N899, N643, N910, N2824, N655, N903, N574, N251, N586, N252, N603, N608, N253, N2815, N2226, N263, N2829, N2214, N266, N2818, N1975, N269, N2821, N1919, N272, N277, N280, N921, N922, N290, N926, N306, n_75, N682, N685, N550, N601, N602, N275, N1344, N1513, N2753, N1267, N1487, N2669, N1352, N1472, N2754, N1433, N2671, N1484, N2755, N1438, N2673, N1150, N1376, N1464, N2756, N1412, N2675, N1232, N1517, N2779, N1489, N2724, N1243, N1358, N2780, N2726, N1249, N2781, N2728, N2782, N2730, N1158, N1748, N2783, N1712, N2732, N1246, N1521, N2762, N1493, N2682, N1478, N1526, N2784, N1434, N1495, N2735, N1370, N1481, N2785, N1439, N2737, N1162, N2786, N1068, N2739, N2787, N2741, N1235, N1364, N2767, N1121, N2688, N1529, N2768, N1498, N2690, N1159, N2232, N1348, N2850, N2857, N991, N2266, N2386, N2279, N1163, N1706, N893, N2024, N1350, N2854, N2861, N896, N2272, N2427, N1167, N1825, N1155, N1496, N1157, N612, N2851, N2858, N2244, N2234, N2863, N2862, N2236, N2230, N2852, N2859, N2026, N2008, N2853, N2860, N1979, N1941, N1171, N1188, N1802, N1858, N1889, N2062, N2078, N2081, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N923, N2384, N2800, N2881, N886, N2882, N887, N2886, N2887, N2888, N2889, N2890, N2899, N1965, N1968, N2773, N2776, N2003, N2897, N1440, N1746, N1809, N1546, N1444, N1769, N1528, N1567, N1532, N1821, N1264, N1459, N1460, N1638, N1510, N1386, N1855, N1561, N1396, N1448, N1346, N1826, N1319, N1795, N1796, N1398, N1759, N1554, N1636, N1530, N1882, N1557, N1458, N1568, N1531, N1772, N1334, N1388, N1454, N1594, N1688, N1576, N2240, N2222, N2876, N2866, N2537, N2540, N2543, N2546, N2549, N2552, N2555, N2594, N2597, N2600, N2603, N2606, n_59, n_66, N2611, N2614, N2617, N2620, n_71, N2385, N1742, N1671, N2041, N2004, N2880, N2870, N2426, N1850, N1527, N2877, N2867, N2256, N2883, N2875, N2361, N2375, N2250, N2878, N2868, N2129, N2143, N2047, N2879, N2869, N2119, N2012, N2558, N2561, N2564, N2567, N2639, N2642, N2645, N2648, N2570, N2573, N2576, N2651, N2655, N2658, N2661, N2664, N1920, N1976, N2005, N2215, N2223, N2227, n_76, n_77, n_78, N2811, N2891, N2871, N2892, N2873, N2827, N2018, N2828, N2019, N2807, N2808, N2809, N2810, N2040, N2898, N2023, N2895, N1774, N1838, N1708, N1784, N1798, N1740, N1596, N1878, N1848, N1723, N1913, N1885, N1884, N1852, N1788, N1720, N1685, N1936, N1911, N1830, N1801, N2253, N2745, n_79, n_80, N2746, n_83, n_86, n_81, n_82, n_84, n_85, N1857, N2353, N2067, N2000, N2036, N1898, N2016, N1571, N2896, N2340, N2104, N2670, N2672, N2674, N2676, N2725, N2727, N2729, N2731, N2683, N2689, N2691, N2733, N2736, N2738, N2740, N2742, N2843, N2846, N1822, N1883, N1915, N1672, N2014, N1910, N1773, N1947, N1912, N1827, N1741, N1987, N1938, N2747, N2750, N2038, N2052, N2020, N2055, N2022, N2872, N2874, N2789, N2060, N2076, N2077;
	wire N2789_key, N2022_key, N1_key, N4_key, N7_key, N10_key, N13_key, N16_key, N19_key, N22_key, N25_key, N28_key, N31_key, N34_key, N37_key, N40_key, N43_key, N46_key, N49_key, N53_key, N56_key, N60_key, N63_key, N66_key, N69_key, N72_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25;
	assign N1160 = ~( N592 & N1_key );
	assign N1443 = ~( N1352 & N1_key );
	assign N2720 = ~( N1_key & N2670 );
	assign N190 = ~N1_key;
	assign N1309 = ~( N197 & N4_key );
	assign N1387 = ~( N1232 & N4_key );
	assign N2721 = ~( N4_key & N2672 );
	assign N194 = ~N4_key;
	assign N1206 = ~( N194 & N7_key );
	assign N1397 = ~( N1243 & N7_key );
	assign N2722 = ~( N7_key & N2674 );
	assign N197 = ~N7_key;
	assign N1054 = ~( N216 & N10_key );
	assign N1226 = ~( N239 & N10_key );
	assign N1345 = ~( N1249 & N10_key );
	assign N2723 = ~( N10_key & N2676 );
	assign N201 = ~N10_key;
	assign N1119 = ~( N216 & N13_key );
	assign N1447 = ~( N1358 & N13_key );
	assign N2757 = ~( N13_key & N2725 );
	assign N206 = ~N13_key;
	assign N1128 = ~( N216 & N16_key );
	assign N1311 = ~( N212 & N16_key );
	assign N2758 = ~( N16_key & N2727 );
	assign N209 = ~N16_key;
	assign N1132 = ~( N225 & N19_key );
	assign N1210 = ~( N209 & N19_key );
	assign N2759 = ~( N19_key & N2729 );
	assign N212 = ~N19_key;
	assign N1055 = ~( N201 & N22_key );
	assign N1120 = ~( N206 & N22_key );
	assign N1129 = ~( N209 & N22_key );
	assign N2760 = ~( N22_key & N2731 );
	assign N216 = ~N22_key;
	assign N1063 = ~( N239 & N25_key );
	assign N1678 = ~( N1521 & N25_key );
	assign N2761 = ~( N25_key & N2733 );
	assign N220 = ~N25_key;
	assign N1130 = ~( N243 & N28_key );
	assign N1133 = ~( N212 & N28_key );
	assign N1453 = ~( N1364 & N28_key );
	assign N2734 = ~( N28_key & N2683 );
	assign N225 = ~N28_key;
	assign N1389 = ~( N1235 & N31_key );
	assign N1457 = ~( N1370 & N31_key );
	assign N2763 = ~( N31_key & N2736 );
	assign N229 = ~N31_key;
	assign N1315 = ~( N235 & N34_key );
	assign N1399 = ~( N1246 & N34_key );
	assign N2764 = ~( N34_key & N2738 );
	assign N232 = ~N34_key;
	assign N1067 = ~( N655 & N37_key );
	assign N1221 = ~( N232 & N37_key );
	assign N2765 = ~( N37_key & N2740 );
	assign N235 = ~N37_key;
	assign N1064 = ~( N220 & N40_key );
	assign N1317 = ~( N201 & N40_key );
	assign N2766 = ~( N40_key & N2742 );
	assign N239 = ~N40_key;
	assign N1122 = ~( N724 & N43_key );
	assign N1131 = ~( N225 & N43_key );
	assign N1313 = ~( N247 & N43_key );
	assign N2743 = ~( N43_key & N2689 );
	assign N243 = ~N43_key;
	assign N1214 = ~( N243 & N46_key );
	assign N1462 = ~( N1158 & N46_key );
	assign N2744 = ~( N46_key & N2691 );
	assign N247 = ~N46_key;
	assign N592 = ( N49_key & N253 & N275 );
	assign N907 = ~( N49_key & N612 );
	assign N2812 = ( N49_key & N612 & N94 & N2789_key );
	assign N724 = ( N53_key & N253 & N275 );
	assign N899 = ~( N53_key & N612 );
	assign N643 = ( N56_key & N69_key & N275 );
	assign N910 = ~( N56_key & N608 );
	assign N2824 = ( N56_key & N608 & N94 & N2789_key );
	assign N655 = ( N60_key & N69_key & N275 );
	assign N903 = ~( N60_key & N608 );
	assign N574 = ( N63_key & N275 );
	assign N251 = ~( N63_key & N88 );
	assign N586 = ( N66_key & N275 );
	assign N252 = ~( N66_key & N91 );
	assign N603 = ~( N69_key & N72_key );
	assign N608 = ~( N69_key & N290 );
	assign N253 = ~N72_key;
	assign N2815 = ( N76 & N94 & N2789_key );
	assign N2226 = ~( N2081 & N76 );
	assign N263 = ~N76;
	assign N2829 = ( N79 & N94 & N2789_key );
	assign N2214 = ~( N2062 & N79 );
	assign N266 = ~N79;
	assign N2818 = ( N82 & N94 & N2789_key );
	assign N1975 = ~( N1858 & N82 );
	assign N269 = ~N82;
	assign N2821 = ( N85 & N94 & N2789_key );
	assign N1919 = ~( N1802 & N85 );
	assign N272 = ~N85;
	assign N277 = ~N88;
	assign N280 = ~N91;
	assign N921 = ~( N277 & N94 & N104 & N603 );
	assign N922 = ~( N280 & N94 & N104 & N603 );
	assign N290 = ~N94;
	assign N926 = ( N99 & N275 & N603 );
	assign N306 = ~N99;
	assign n_75 = ( N275 & N2279 & N99 & N2747 );
	assign N682 = ( N251 & N104 );
	assign N685 = ( N252 & N104 );
	assign N550 = ~( N306 & N104 );
	assign N601 = ~( N104 & N277 );
	assign N602 = ~( N104 & N280 );
	assign N275 = ~N104;
	assign N1344 = ~( N1267 & N1160 );
	assign N1513 = ~( N1443 & N1487 );
	assign N2753 = ~( N2669 & N2720 );
	assign N1267 = ~( N190 & N1159 );
	assign N1487 = ~( N190 & N1444 );
	assign N2669 = ~( N2558 & N190 );
	assign N1352 = ~( N1309 & N1206 );
	assign N1472 = ~( N1387 & N1433 );
	assign N2754 = ~( N2671 & N2721 );
	assign N1433 = ~( N194 & N1386 );
	assign N2671 = ~( N2561 & N194 );
	assign N1484 = ~( N1397 & N1438 );
	assign N2755 = ~( N2673 & N2722 );
	assign N1438 = ~( N197 & N1396 );
	assign N2673 = ~( N2564 & N197 );
	assign N1150 = ~( N1054 & N1055 );
	assign N1376 = ~( N1317 & N1226 );
	assign N1464 = ~( N1345 & N1412 );
	assign N2756 = ~( N2675 & N2723 );
	assign N1412 = ~( N201 & N1346 );
	assign N2675 = ~( N2567 & N201 );
	assign N1232 = ~( N1119 & N1120 );
	assign N1517 = ~( N1447 & N1489 );
	assign N2779 = ~( N2724 & N2757 );
	assign N1489 = ~( N206 & N1448 );
	assign N2724 = ~( N2639 & N206 );
	assign N1243 = ~( N1128 & N1129 );
	assign N1358 = ~( N1311 & N1210 );
	assign N2780 = ~( N2726 & N2758 );
	assign N2726 = ~( N2642 & N209 );
	assign N1249 = ~( N1132 & N1133 );
	assign N2781 = ~( N2728 & N2759 );
	assign N2728 = ~( N2645 & N212 );
	assign N2782 = ~( N2730 & N2760 );
	assign N2730 = ~( N2648 & N216 );
	assign N1158 = ~( N1063 & N1064 );
	assign N1748 = ~( N1678 & N1712 );
	assign N2783 = ~( N2732 & N2761 );
	assign N1712 = ~( N220 & N1554 );
	assign N2732 = ~( N2651 & N220 );
	assign N1246 = ~( N1130 & N1131 );
	assign N1521 = ~( N1453 & N1493 );
	assign N2762 = ~( N2682 & N2734 );
	assign N1493 = ~( N225 & N1454 );
	assign N2682 = ~( N2570 & N225 );
	assign N1478 = ~( N1389 & N1434 );
	assign N1526 = ~( N1457 & N1495 );
	assign N2784 = ~( N2735 & N2763 );
	assign N1434 = ~( N229 & N1388 );
	assign N1495 = ~( N229 & N1458 );
	assign N2735 = ~( N2655 & N229 );
	assign N1370 = ~( N1315 & N1221 );
	assign N1481 = ~( N1399 & N1439 );
	assign N2785 = ~( N2737 & N2764 );
	assign N1439 = ~( N232 & N1398 );
	assign N2737 = ~( N2658 & N232 );
	assign N1162 = ~( N1067 & N1068 );
	assign N2786 = ~( N2739 & N2765 );
	assign N1068 = ~( N235 & N896 );
	assign N2739 = ~( N2661 & N235 );
	assign N2787 = ~( N2741 & N2766 );
	assign N2741 = ~( N2664 & N239 );
	assign N1235 = ~( N1121 & N1122 );
	assign N1364 = ~( N1313 & N1214 );
	assign N2767 = ~( N2688 & N2743 );
	assign N1121 = ~( N243 & N991 );
	assign N2688 = ~( N2573 & N243 );
	assign N1529 = ~( N1462 & N1498 );
	assign N2768 = ~( N2690 & N2744 );
	assign N1498 = ~( N247 & N1319 );
	assign N2690 = ~( N2576 & N247 );
	assign N1159 = ~N592;
	assign N2232 = ~( N907 & N2223 );
	assign N1348 = ~N907;
	assign N2850 = ~( N2812 & N2076 );
	assign N2857 = ~N2812;
	assign N991 = ~N724;
	assign N2266 = ( N899 & N2240 );
	assign N2386 = ( N899 & N2253 );
	assign N2279 = ~( N2067 & N2012 & N2047 & N2250 & N899 & N2256 & N2253 & N903 );
	assign N1163 = ~N899;
	assign N1706 = ~( N643 & N1672 );
	assign N893 = ~N643;
	assign N2024 = ~( N910 & N2005 );
	assign N1350 = ~N910;
	assign N2854 = ~( N2824 & N1938 );
	assign N2861 = ~N2824;
	assign N896 = ~N655;
	assign N2272 = ( N903 & N2244 );
	assign N2427 = ( N903 & N2256 );
	assign N1167 = ~N903;
	assign N1825 = ~( N574 & N1796 );
	assign N1155 = ~N574;
	assign N1496 = ~( N586 & N1460 );
	assign N1157 = ~N586;
	assign N612 = ~( N253 & N290 );
	assign N2851 = ~( N2815 & N2077 );
	assign N2858 = ~N2815;
	assign N2244 = ~( N2226 & N2234 );
	assign N2234 = ~( N263 & N2227 );
	assign N2863 = ~( N2829 & N1947 );
	assign N2862 = ~N2829;
	assign N2236 = ~( N2214 & N2230 );
	assign N2230 = ~( N266 & N2215 );
	assign N2852 = ~( N2818 & N1915 );
	assign N2859 = ~N2818;
	assign N2026 = ~( N1975 & N2008 );
	assign N2008 = ~( N269 & N1976 );
	assign N2853 = ~( N2821 & N1857 );
	assign N2860 = ~N2821;
	assign N1979 = ~( N1919 & N1941 );
	assign N1941 = ~( N272 & N1920 );
	assign N1171 = ~( N921 & N923 );
	assign N1188 = ~( N922 & N923 );
	assign N1802 = ~( N1742 & N290 );
	assign N1858 = ~( N1798 & N290 );
	assign N1889 = ~( N1830 & N290 );
	assign N2062 = ~( N2040 & N290 );
	assign N2078 = ~( N2060 & N290 );
	assign N2081 = ~( N2055 & N290 );
	assign N2627 = ~( N2266 & N2427 & N2340 & N2104 & N926 );
	assign N2628 = ~( N2386 & N2272 & N2340 & N2104 & N926 );
	assign N2629 = ~( N2386 & N2427 & N2361 & N2104 & N926 );
	assign N2630 = ~( N2386 & N2427 & N2340 & N2129 & N926 );
	assign N2631 = ~( N2386 & N2427 & N2340 & N2119 & N926 );
	assign N2632 = ~( N2386 & N2427 & N2353 & N2104 & N926 );
	assign N2633 = ~( N2386 & N2426 & N2340 & N2104 & N926 );
	assign N2634 = ~( N2385 & N2427 & N2340 & N2104 & N926 );
	assign N923 = ~N926;
	assign N2384 = ( N275 & N2279 & N306 );
	assign N2800 = ( n_75 & n_76 & n_77 & n_78 );
	assign N2881 = ~( N682 & N2872 );
	assign N886 = ~N682;
	assign N2882 = ~( N685 & N2874 );
	assign N887 = ~N685;
	assign N2886 = ( N2876 & N550 );
	assign N2887 = ( N550 & N2877 );
	assign N2888 = ( N550 & N2878 );
	assign N2889 = ( N2879 & N550 );
	assign N2890 = ( N550 & N2880 );
	assign N2899 = ( N2898 & N550 );
	assign N1965 = ( N1910 & N601 );
	assign N1968 = ( N602 & N1912 );
	assign N2773 = ( N2745 & N275 );
	assign N2776 = ( N2746 & N275 );
	assign N2003 = ~( N1947 & N1344 );
	assign N2897 = ~( N1344 & N2896 );
	assign N1440 = ~N1344;
	assign N1746 = ~( N1517 & N1513 );
	assign N1809 = ~( N1513 & N1521 );
	assign N1546 = ~N1513;
	assign N1444 = ~N1352;
	assign N1769 = ~( N1472 & N1741 );
	assign N1528 = ~N1472;
	assign N1567 = ~( N1484 & N1531 );
	assign N1532 = ~N1484;
	assign N1821 = ~( N1774 & N1150 );
	assign N1264 = ~N1150;
	assign N1459 = ~( N1376 & N1157 );
	assign N1460 = ~N1376;
	assign N1638 = ~( N1576 & N1464 );
	assign N1510 = ~N1464;
	assign N1386 = ~N1232;
	assign N1855 = ~( N1788 & N1517 );
	assign N1561 = ~N1517;
	assign N1396 = ~N1243;
	assign N1448 = ~N1358;
	assign N1346 = ~N1249;
	assign N1826 = ~( N1788 & N1158 );
	assign N1319 = ~N1158;
	assign N1795 = ~( N1748 & N1155 );
	assign N1796 = ~N1748;
	assign N1398 = ~N1246;
	assign N1759 = ~( N1526 & N1521 );
	assign N1554 = ~N1521;
	assign N1636 = ~( N1478 & N1576 );
	assign N1530 = ~N1478;
	assign N1882 = ~( N1838 & N1526 );
	assign N1557 = ~N1526;
	assign N1458 = ~N1370;
	assign N1568 = ~( N1481 & N1532 );
	assign N1531 = ~N1481;
	assign N1772 = ~( N1723 & N1162 );
	assign N1334 = ~N1162;
	assign N1388 = ~N1235;
	assign N1454 = ~N1364;
	assign N1594 = ~( N1529 & N1530 );
	assign N1688 = ~( N1510 & N1529 );
	assign N1576 = ~N1529;
	assign N2240 = ~( N2222 & N2232 );
	assign N2222 = ~( N2078 & N1348 );
	assign N2876 = ~( N2866 & N2850 );
	assign N2866 = ~( N2052 & N2857 );
	assign N2537 = ~( N2266 & N2272 & N2361 & N2104 & N1171 );
	assign N2540 = ~( N2266 & N2272 & N2340 & N2129 & N1171 );
	assign N2543 = ~( N2266 & N2272 & N2340 & N2119 & N1171 );
	assign N2546 = ~( N2266 & N2272 & N2353 & N2104 & N1171 );
	assign N2549 = ~( N2266 & N2272 & N2375 & N2119 & N1188 );
	assign N2552 = ~( N2266 & N2272 & N2361 & N2143 & N1188 );
	assign N2555 = ~( N2266 & N2272 & N2375 & N2129 & N1188 );
	assign N2594 = ~( N2266 & N2427 & N2361 & N2129 & N1171 );
	assign N2597 = ~( N2266 & N2427 & N2361 & N2119 & N1171 );
	assign N2600 = ~( N2266 & N2427 & N2375 & N2104 & N1171 );
	assign N2603 = ~( N2266 & N2427 & N2340 & N2143 & N1171 );
	assign N2606 = ~( N2266 & N2427 & N2353 & N2129 & N1188 );
	assign n_59 = ( N2266 & N2272 );
	assign n_66 = ( N2266 & N2427 );
	assign N2611 = ~( N2386 & N2272 & N2361 & N2129 & N1188 );
	assign N2614 = ~( N2386 & N2272 & N2361 & N2119 & N1188 );
	assign N2617 = ~( N2386 & N2272 & N2375 & N2104 & N1188 );
	assign N2620 = ~( N2386 & N2272 & N2353 & N2129 & N1188 );
	assign n_71 = ( N2386 & N2272 );
	assign N2385 = ( N1163 & N2253 );
	assign N1742 = ~( N1671 & N1706 );
	assign N1671 = ~( N1596 & N893 );
	assign N2041 = ~( N2004 & N2024 );
	assign N2004 = ~( N1889 & N1350 );
	assign N2880 = ~( N2870 & N2854 );
	assign N2870 = ~( N1830 & N2861 );
	assign N2426 = ( N1167 & N2256 );
	assign N1850 = ~( N1795 & N1825 );
	assign N1527 = ~( N1459 & N1496 );
	assign N2877 = ~( N2867 & N2851 );
	assign N2867 = ~( N2055 & N2858 );
	assign N2256 = ~N2244;
	assign N2883 = ~( N2875 & N2863 );
	assign N2875 = ~( N1913 & N2862 );
	assign N2361 = ( N2067 & N2236 );
	assign N2375 = ( N2041 & N2236 );
	assign N2250 = ~N2236;
	assign N2878 = ~( N2868 & N2852 );
	assign N2868 = ~( N1798 & N2859 );
	assign N2129 = ( N2012 & N2026 );
	assign N2143 = ( N1979 & N2026 );
	assign N2047 = ~N2026;
	assign N2879 = ~( N2869 & N2853 );
	assign N2869 = ~( N1742 & N2860 );
	assign N2119 = ( N1979 & N2047 );
	assign N2012 = ~N1979;
	assign N2558 = ( N2361 & N2104 & N1171 & n_59 );
	assign N2561 = ( N2340 & N2129 & N1171 & n_59 );
	assign N2564 = ( N2340 & N2119 & N1171 & n_59 );
	assign N2567 = ( N2353 & N2104 & N1171 & n_59 );
	assign N2639 = ( N2361 & N2129 & N1171 & n_66 );
	assign N2642 = ( N2361 & N2119 & N1171 & n_66 );
	assign N2645 = ( N2375 & N2104 & N1171 & n_66 );
	assign N2648 = ( N2340 & N2143 & N1171 & n_66 );
	assign N2570 = ( N2375 & N2119 & N1188 & n_59 );
	assign N2573 = ( N2361 & N2143 & N1188 & n_59 );
	assign N2576 = ( N2375 & N2129 & N1188 & n_59 );
	assign N2651 = ( N2353 & N2129 & N1188 & n_66 );
	assign N2655 = ( N2361 & N2129 & N1188 & n_71 );
	assign N2658 = ( N2361 & N2119 & N1188 & n_71 );
	assign N2661 = ( N2375 & N2104 & N1188 & n_71 );
	assign N2664 = ( N2353 & N2129 & N1188 & n_71 );
	assign N1920 = ~N1802;
	assign N1976 = ~N1858;
	assign N2005 = ~N1889;
	assign N2215 = ~N2062;
	assign N2223 = ~N2078;
	assign N2227 = ~N2081;
	assign n_76 = ( N2750 & N2627 & N2628 );
	assign n_77 = ( N2629 & N2630 & N2631 );
	assign n_78 = ( N2632 & N2633 & N2634 );
	assign N2811 = ~( N2384 | N2800 );
	assign N2891 = ~( N2871 & N2881 );
	assign N2871 = ~( N2843 & N886 );
	assign N2892 = ~( N2873 & N2882 );
	assign N2873 = ~( N2846 & N887 );
	assign N2827 = ~( N1965 & N2808 );
	assign N2018 = ~N1965;
	assign N2828 = ~( N1968 & N2810 );
	assign N2019 = ~N1968;
	assign N2807 = ~( N2773 & N2018 );
	assign N2808 = ~N2773;
	assign N2809 = ~( N2776 & N2019 );
	assign N2810 = ~N2776;
	assign N2040 = ~( N2023 & N2003 );
	assign N2898 = ~( N2895 & N2897 );
	assign N2023 = ~( N1440 & N1913 );
	assign N2895 = ~( N2883 & N1440 );
	assign N1774 = ~( N1708 & N1746 );
	assign N1838 = ~( N1809 & N1784 );
	assign N1708 = ~( N1546 & N1561 );
	assign N1784 = ~( N1554 & N1546 );
	assign N1798 = ~( N1740 & N1769 );
	assign N1740 = ~( N1685 & N1528 );
	assign N1596 = ~( N1567 & N1568 );
	assign N1878 = ~( N1821 & N1848 );
	assign N1848 = ~( N1264 & N1822 );
	assign N1723 = ~( N1638 & N1688 );
	assign N1913 = ~( N1855 & N1885 );
	assign N1885 = ~( N1561 & N1827 );
	assign N1884 = ~( N1826 & N1852 );
	assign N1852 = ~( N1319 & N1827 );
	assign N1788 = ~( N1720 & N1759 );
	assign N1720 = ~( N1554 & N1557 );
	assign N1685 = ~( N1594 & N1636 );
	assign N1936 = ~( N1882 & N1911 );
	assign N1911 = ~( N1557 & N1883 );
	assign N1830 = ~( N1772 & N1801 );
	assign N1801 = ~( N1334 & N1773 );
	assign N2253 = ~N2240;
	assign N2745 = ~( N2537 & N2540 & N2543 & N2546 & N2594 & N2597 & N2600 & N2603 );
	assign n_79 = ( N2537 & N2540 );
	assign n_80 = ( N2543 & N2546 );
	assign N2746 = ~( N2606 & N2549 & N2611 & N2614 & N2617 & N2620 & N2552 & N2555 );
	assign n_83 = ( N2606 & N2549 );
	assign n_86 = ( N2552 & N2555 );
	assign n_81 = ( N2594 & N2597 );
	assign n_82 = ( N2600 & N2603 );
	assign n_84 = ( N2611 & N2614 );
	assign n_85 = ( N2617 & N2620 );
	assign N1857 = ~N1742;
	assign N2353 = ( N2041 & N2250 );
	assign N2067 = ~N2041;
	assign N2000 = ~( N1878 & N1850 );
	assign N2036 = ~( N1850 & N1910 );
	assign N1898 = ~N1850;
	assign N2016 = ~( N1936 & N1527 );
	assign N1571 = ~N1527;
	assign N2896 = ~N2883;
	assign N2340 = ( N2067 & N2250 );
	assign N2104 = ( N2012 & N2047 );
	assign N2670 = ~N2558;
	assign N2672 = ~N2561;
	assign N2674 = ~N2564;
	assign N2676 = ~N2567;
	assign N2725 = ~N2639;
	assign N2727 = ~N2642;
	assign N2729 = ~N2645;
	assign N2731 = ~N2648;
	assign N2683 = ~N2570;
	assign N2689 = ~N2573;
	assign N2691 = ~N2576;
	assign N2733 = ~N2651;
	assign N2736 = ~N2655;
	assign N2738 = ~N2658;
	assign N2740 = ~N2661;
	assign N2742 = ~N2664;
	assign N2843 = ~( N2807 & N2827 );
	assign N2846 = ~( N2809 & N2828 );
	assign N1822 = ~N1774;
	assign N1883 = ~N1838;
	assign N1915 = ~N1798;
	assign N1672 = ~N1596;
	assign N2014 = ~( N1878 & N1898 );
	assign N1910 = ~N1878;
	assign N1773 = ~N1723;
	assign N1947 = ~N1913;
	assign N1912 = ~N1884;
	assign N1827 = ~N1788;
	assign N1741 = ~N1685;
	assign N1987 = ~N1936;
	assign N1938 = ~N1830;
	assign N2747 = ( n_79 & n_80 & n_81 & n_82 );
	assign N2750 = ( n_83 & n_84 & n_85 & n_86 );
	assign N2038 = ~( N2020 & N2000 );
	assign N2052 = ~( N2036 & N2014 );
	assign N2020 = ~( N1898 & N1910 );
	assign N2055 = ~( N2022_key & N2016 );
	assign N2022 = ~( N1987 & N1571 );
	assign N2872 = ~N2843;
	assign N2874 = ~N2846;
	assign N2789 = ~( N2747 & N2750 );
	assign N2060 = ~N2038;
	assign N2076 = ~N2052;
	assign N2077 = ~N2055;
	assign N2789_key = ~( N2789 ^ key_0 );
	assign N2022_key = ~( N2022 ^ key_1 );
	assign N1_key = ~( N1 ^ key_2 );
	assign N4_key = ~( N4 ^ key_3 );
	assign N7_key = ~( N7 ^ key_4 );
	assign N10_key = ~( N10 ^ key_5 );
	assign N13_key = ~( N13 ^ key_6 );
	assign N16_key = ~( N16 ^ key_7 );
	assign N19_key = ~( N19 ^ key_8 );
	assign N22_key = ~( N22 ^ key_9 );
	assign N25_key = ~( N25 ^ key_10 );
	assign N28_key = ~( N28 ^ key_11 );
	assign N31_key = ~( N31 ^ key_12 );
	assign N34_key = ~( N34 ^ key_13 );
	assign N37_key = ~( N37 ^ key_14 );
	assign N40_key = ~( N40 ^ key_15 );
	assign N43_key = ~( N43 ^ key_16 );
	assign N46_key = ~( N46 ^ key_17 );
	assign N49_key = ~( N49 ^ key_18 );
	assign N53_key = ~( N53 ^ key_19 );
	assign N56_key = ~( N56 ^ key_20 );
	assign N60_key = ~( N60 ^ key_21 );
	assign N63_key = ~( N63 ^ key_22 );
	assign N66_key = ~( N66 ^ key_23 );
	assign N69_key = ~( N69 ^ key_24 );
	assign N72_key = ~( N72 ^ key_25 );
endmodule
