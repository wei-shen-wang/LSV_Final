module c1355(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355);
	input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29;
	output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
	wire G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, G266, G314, G362, G394, G1132, G1228, G278, G323, G371, G400, G1159, G1246, G281, G329, G372, G404, G1162, G1248, G335, G373, G408, G1165, G1250, G284, G317, G374, G397, G1168, G1252, G375, G401, G1171, G1254, G287, G376, G405, G1174, G1256, G377, G409, G1177, G1258, G290, G338, G378, G410, G1180, G1260, G344, G379, G414, G1183, G1262, G293, G350, G380, G418, G1186, G1264, G320, G363, G398, G1135, G1230, G356, G381, G422, G1189, G1266, G296, G382, G411, G1192, G1268, G383, G415, G1195, G1270, G299, G384, G419, G1198, G1272, G385, G423, G1201, G1274, G302, G341, G386, G412, G1204, G1276, G347, G387, G416, G1207, G1278, G305, G353, G388, G420, G1210, G1280, G359, G389, G424, G1213, G1282, G308, G390, G413, G1216, G1284, G269, G326, G364, G402, G1138, G1232, G391, G417, G1219, G1286, G311, G392, G421, G1222, G1288, G393, G425, G1225, G1290, G242, G245, G248, G251, G254, G257, G260, G332, G365, G406, G1141, G1234, G263, G272, G366, G395, G1144, G1236, G367, G399, G1147, G1238, G275, G368, G403, G1150, G1240, G369, G407, G1153, G1242, G370, G396, G1156, G1244, G426, G474, G1229, G1292, G438, G483, G1247, G1301, G441, G489, G1249, G1302, G495, G1251, G1303, G444, G477, G1253, G1304, G1255, G1305, G447, G1257, G1306, G1259, G1307, G450, G498, G1261, G1308, G504, G1263, G1309, G453, G510, G1265, G1310, G480, G1231, G1293, G516, G1267, G1311, G456, G1269, G1312, G1271, G1313, G459, G1273, G1314, G1275, G1315, G462, G501, G1277, G1316, G507, G1279, G1317, G465, G513, G1281, G1318, G519, G1283, G1319, G468, G1285, G1320, G429, G486, G1233, G1294, G1287, G1321, G471, G1289, G1322, G1291, G1323, G730, G754, G733, G756, G736, G758, G739, G760, G742, G762, G745, G764, G748, G766, G492, G1235, G1295, G751, G768, G432, G1237, G1296, G1239, G1297, G435, G1241, G1298, G1243, G1299, G1245, G1300, G522, G570, G546, G586, G1324, G528, G574, G549, G589, G1333, G575, G552, G591, G1334, G555, G593, G1335, G531, G576, G587, G1336, G1337, G577, G1338, G1339, G534, G578, G558, G594, G1340, G561, G596, G1341, G579, G564, G598, G1342, G588, G1325, G567, G600, G1343, G537, G580, G1344, G1345, G581, G1346, G1347, G540, G582, G595, G1348, G597, G1349, G583, G599, G1350, G601, G1351, G543, G584, G1352, G571, G590, G1326, G1353, G585, G1354, G1355, G755, G770, G757, G773, G759, G776, G761, G779, G763, G782, G765, G785, G767, G788, G592, G1327, G769, G791, G525, G572, G1328, G1329, G573, G1330, G1331, G1332, G602, G642, G612, G645, G648, G651, G617, G622, G654, G657, G660, G663, G627, G632, G637, G794, G819, G797, G821, G800, G823, G803, G825, G806, G827, G809, G829, G812, G831, G815, G833, G607, G666, G672, G690, G694, G818, G669, G692, G695, G820, G822, G824, G675, G693, G697, G678, G684, G698, G702, G826, G828, G830, G832, G687, G699, G704, G681, G700, G703, G701, G705, G834, G847, G860, G873, G925, G886, G912, G899, G691, G696, G706, G712, G709, G715, G718, G724, G727, G721, G1036, G1048, G1060, G1072, AND4_3_inw1, G938, n_78, G1039, G1051, G1063, G1075, AND4_2_inw1, G939, n_80, G1042, G1054, G1066, G1078, AND4_1_inw2, G940, g10_inw1, g14_inw1, G1045, G1057, G1069, G1081, AND4_0_inw2, G943, g12_inw1, g16_inw1, G1084, G1096, G1108, G1120, AND4_7_inw1, G954, n_74, G1087, G1099, G1111, G1123, AND4_6_inw1, G950, n_76, G1090, G1102, G1114, G1126, AND4_5_inw2, G953, g2_inw1, g6_inw1, G1093, G1105, G1117, G1129, AND4_4_inw2, G951, g4_inw1, g8_inw1, G981, AND4_0_inw1, AND4_1_inw1, g10_inw2, g12_inw2, G980, g14_inw2, g16_inw2, G979, AND4_2_inw2, AND4_3_inw2, G1016, G1026, G978, G1021, G1031, G985, AND4_4_inw1, AND4_5_inw1, g2_inw2, g4_inw2, G984, g6_inw2, g8_inw2, G983, AND4_6_inw2, AND4_7_inw2, G996, G1006, G982, G1001, G1011, OR4_0_inw2, OR4_0_inw1, OR4_1_inw2, OR4_1_inw1, G986, G991;
	wire G991_key, G986_key, OR4_1_inw1_key, AND4_7_inw1_key, AND4_6_inw1_key, AND4_5_inw2_key, AND4_4_inw2_key, G985_key, AND4_4_inw1_key, AND4_5_inw1_key, G984_key, G983_key, AND4_6_inw2_key, AND4_7_inw2_key, G982_key, OR4_1_inw2_key, AND4_3_inw1_key, AND4_2_inw1_key, AND4_1_inw2_key, AND4_0_inw2_key, G981_key, AND4_0_inw1_key, AND4_1_inw1_key, G980_key, G979_key, AND4_2_inw2_key, AND4_3_inw2_key, G978_key, OR4_0_inw2_key, OR4_0_inw1_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29;
	assign G266 = ~( G1 & G2 );
	assign G314 = ~( G1 & G5 );
	assign G362 = ~( G1 & G266 );
	assign G394 = ~( G1 & G314 );
	assign G1132 = ~( G1 & G1036 );
	assign G1228 = ~( G1 & G1132 );
	assign G278 = ~( G9 & G10 );
	assign G323 = ~( G10 & G14 );
	assign G371 = ~( G10 & G278 );
	assign G400 = ~( G10 & G323 );
	assign G1159 = ~( G10 & G1063 );
	assign G1246 = ~( G10 & G1159 );
	assign G281 = ~( G11 & G12 );
	assign G329 = ~( G11 & G15 );
	assign G372 = ~( G11 & G281 );
	assign G404 = ~( G11 & G329 );
	assign G1162 = ~( G11 & G1066 );
	assign G1248 = ~( G11 & G1162 );
	assign G335 = ~( G12 & G16 );
	assign G373 = ~( G12 & G281 );
	assign G408 = ~( G12 & G335 );
	assign G1165 = ~( G12 & G1069 );
	assign G1250 = ~( G12 & G1165 );
	assign G284 = ~( G13 & G14 );
	assign G317 = ~( G9 & G13 );
	assign G374 = ~( G13 & G284 );
	assign G397 = ~( G13 & G317 );
	assign G1168 = ~( G13 & G1072 );
	assign G1252 = ~( G13 & G1168 );
	assign G375 = ~( G14 & G284 );
	assign G401 = ~( G14 & G323 );
	assign G1171 = ~( G14 & G1075 );
	assign G1254 = ~( G14 & G1171 );
	assign G287 = ~( G15 & G16 );
	assign G376 = ~( G15 & G287 );
	assign G405 = ~( G15 & G329 );
	assign G1174 = ~( G15 & G1078 );
	assign G1256 = ~( G15 & G1174 );
	assign G377 = ~( G16 & G287 );
	assign G409 = ~( G16 & G335 );
	assign G1177 = ~( G16 & G1081 );
	assign G1258 = ~( G16 & G1177 );
	assign G290 = ~( G17 & G18 );
	assign G338 = ~( G17 & G21 );
	assign G378 = ~( G17 & G290 );
	assign G410 = ~( G17 & G338 );
	assign G1180 = ~( G17 & G1084 );
	assign G1260 = ~( G17 & G1180 );
	assign G344 = ~( G18 & G22 );
	assign G379 = ~( G18 & G290 );
	assign G414 = ~( G18 & G344 );
	assign G1183 = ~( G18 & G1087 );
	assign G1262 = ~( G18 & G1183 );
	assign G293 = ~( G19 & G20 );
	assign G350 = ~( G19 & G23 );
	assign G380 = ~( G19 & G293 );
	assign G418 = ~( G19 & G350 );
	assign G1186 = ~( G19 & G1090 );
	assign G1264 = ~( G19 & G1186 );
	assign G320 = ~( G2 & G6 );
	assign G363 = ~( G2 & G266 );
	assign G398 = ~( G2 & G320 );
	assign G1135 = ~( G2 & G1039 );
	assign G1230 = ~( G2 & G1135 );
	assign G356 = ~( G20 & G24 );
	assign G381 = ~( G20 & G293 );
	assign G422 = ~( G20 & G356 );
	assign G1189 = ~( G20 & G1093 );
	assign G1266 = ~( G20 & G1189 );
	assign G296 = ~( G21 & G22 );
	assign G382 = ~( G21 & G296 );
	assign G411 = ~( G21 & G338 );
	assign G1192 = ~( G21 & G1096 );
	assign G1268 = ~( G21 & G1192 );
	assign G383 = ~( G22 & G296 );
	assign G415 = ~( G22 & G344 );
	assign G1195 = ~( G22 & G1099 );
	assign G1270 = ~( G22 & G1195 );
	assign G299 = ~( G23 & G24 );
	assign G384 = ~( G23 & G299 );
	assign G419 = ~( G23 & G350 );
	assign G1198 = ~( G23 & G1102 );
	assign G1272 = ~( G23 & G1198 );
	assign G385 = ~( G24 & G299 );
	assign G423 = ~( G24 & G356 );
	assign G1201 = ~( G24 & G1105 );
	assign G1274 = ~( G24 & G1201 );
	assign G302 = ~( G25 & G26 );
	assign G341 = ~( G25 & G29 );
	assign G386 = ~( G25 & G302 );
	assign G412 = ~( G25 & G341 );
	assign G1204 = ~( G25 & G1108 );
	assign G1276 = ~( G25 & G1204 );
	assign G347 = ~( G26 & G30 );
	assign G387 = ~( G26 & G302 );
	assign G416 = ~( G26 & G347 );
	assign G1207 = ~( G26 & G1111 );
	assign G1278 = ~( G26 & G1207 );
	assign G305 = ~( G27 & G28 );
	assign G353 = ~( G27 & G31 );
	assign G388 = ~( G27 & G305 );
	assign G420 = ~( G27 & G353 );
	assign G1210 = ~( G27 & G1114 );
	assign G1280 = ~( G27 & G1210 );
	assign G359 = ~( G28 & G32 );
	assign G389 = ~( G28 & G305 );
	assign G424 = ~( G28 & G359 );
	assign G1213 = ~( G28 & G1117 );
	assign G1282 = ~( G28 & G1213 );
	assign G308 = ~( G29 & G30 );
	assign G390 = ~( G29 & G308 );
	assign G413 = ~( G29 & G341 );
	assign G1216 = ~( G29 & G1120 );
	assign G1284 = ~( G29 & G1216 );
	assign G269 = ~( G3 & G4 );
	assign G326 = ~( G3 & G7 );
	assign G364 = ~( G3 & G269 );
	assign G402 = ~( G3 & G326 );
	assign G1138 = ~( G3 & G1042 );
	assign G1232 = ~( G3 & G1138 );
	assign G391 = ~( G30 & G308 );
	assign G417 = ~( G30 & G347 );
	assign G1219 = ~( G30 & G1123 );
	assign G1286 = ~( G30 & G1219 );
	assign G311 = ~( G31 & G32 );
	assign G392 = ~( G31 & G311 );
	assign G421 = ~( G31 & G353 );
	assign G1222 = ~( G31 & G1126 );
	assign G1288 = ~( G31 & G1222 );
	assign G393 = ~( G32 & G311 );
	assign G425 = ~( G32 & G359 );
	assign G1225 = ~( G32 & G1129 );
	assign G1290 = ~( G32 & G1225 );
	assign G242 = ( G33 & G41 );
	assign G245 = ( G34 & G41 );
	assign G248 = ( G35 & G41 );
	assign G251 = ( G36 & G41 );
	assign G254 = ( G37 & G41 );
	assign G257 = ( G38 & G41 );
	assign G260 = ( G39 & G41 );
	assign G332 = ~( G4 & G8 );
	assign G365 = ~( G4 & G269 );
	assign G406 = ~( G4 & G332 );
	assign G1141 = ~( G4 & G1045 );
	assign G1234 = ~( G4 & G1141 );
	assign G263 = ( G40 & G41 );
	assign G272 = ~( G5 & G6 );
	assign G366 = ~( G5 & G272 );
	assign G395 = ~( G5 & G314 );
	assign G1144 = ~( G5 & G1048 );
	assign G1236 = ~( G5 & G1144 );
	assign G367 = ~( G6 & G272 );
	assign G399 = ~( G6 & G320 );
	assign G1147 = ~( G6 & G1051 );
	assign G1238 = ~( G6 & G1147 );
	assign G275 = ~( G7 & G8 );
	assign G368 = ~( G7 & G275 );
	assign G403 = ~( G7 & G326 );
	assign G1150 = ~( G7 & G1054 );
	assign G1240 = ~( G7 & G1150 );
	assign G369 = ~( G8 & G275 );
	assign G407 = ~( G8 & G332 );
	assign G1153 = ~( G8 & G1057 );
	assign G1242 = ~( G8 & G1153 );
	assign G370 = ~( G9 & G278 );
	assign G396 = ~( G9 & G317 );
	assign G1156 = ~( G9 & G1060 );
	assign G1244 = ~( G9 & G1156 );
	assign G426 = ~( G362 & G363 );
	assign G474 = ~( G394 & G395 );
	assign G1229 = ~( G1036 & G1132 );
	assign G1292 = ~( G1228 & G1229 );
	assign G438 = ~( G370 & G371 );
	assign G483 = ~( G400 & G401 );
	assign G1247 = ~( G1063 & G1159 );
	assign G1301 = ~( G1246 & G1247 );
	assign G441 = ~( G372 & G373 );
	assign G489 = ~( G404 & G405 );
	assign G1249 = ~( G1066 & G1162 );
	assign G1302 = ~( G1248 & G1249 );
	assign G495 = ~( G408 & G409 );
	assign G1251 = ~( G1069 & G1165 );
	assign G1303 = ~( G1250 & G1251 );
	assign G444 = ~( G374 & G375 );
	assign G477 = ~( G396 & G397 );
	assign G1253 = ~( G1072 & G1168 );
	assign G1304 = ~( G1252 & G1253 );
	assign G1255 = ~( G1075 & G1171 );
	assign G1305 = ~( G1254 & G1255 );
	assign G447 = ~( G376 & G377 );
	assign G1257 = ~( G1078 & G1174 );
	assign G1306 = ~( G1256 & G1257 );
	assign G1259 = ~( G1081 & G1177 );
	assign G1307 = ~( G1258 & G1259 );
	assign G450 = ~( G378 & G379 );
	assign G498 = ~( G410 & G411 );
	assign G1261 = ~( G1084 & G1180 );
	assign G1308 = ~( G1260 & G1261 );
	assign G504 = ~( G414 & G415 );
	assign G1263 = ~( G1087 & G1183 );
	assign G1309 = ~( G1262 & G1263 );
	assign G453 = ~( G380 & G381 );
	assign G510 = ~( G418 & G419 );
	assign G1265 = ~( G1090 & G1186 );
	assign G1310 = ~( G1264 & G1265 );
	assign G480 = ~( G398 & G399 );
	assign G1231 = ~( G1039 & G1135 );
	assign G1293 = ~( G1230 & G1231 );
	assign G516 = ~( G422 & G423 );
	assign G1267 = ~( G1093 & G1189 );
	assign G1311 = ~( G1266 & G1267 );
	assign G456 = ~( G382 & G383 );
	assign G1269 = ~( G1096 & G1192 );
	assign G1312 = ~( G1268 & G1269 );
	assign G1271 = ~( G1099 & G1195 );
	assign G1313 = ~( G1270 & G1271 );
	assign G459 = ~( G384 & G385 );
	assign G1273 = ~( G1102 & G1198 );
	assign G1314 = ~( G1272 & G1273 );
	assign G1275 = ~( G1105 & G1201 );
	assign G1315 = ~( G1274 & G1275 );
	assign G462 = ~( G386 & G387 );
	assign G501 = ~( G412 & G413 );
	assign G1277 = ~( G1108 & G1204 );
	assign G1316 = ~( G1276 & G1277 );
	assign G507 = ~( G416 & G417 );
	assign G1279 = ~( G1111 & G1207 );
	assign G1317 = ~( G1278 & G1279 );
	assign G465 = ~( G388 & G389 );
	assign G513 = ~( G420 & G421 );
	assign G1281 = ~( G1114 & G1210 );
	assign G1318 = ~( G1280 & G1281 );
	assign G519 = ~( G424 & G425 );
	assign G1283 = ~( G1117 & G1213 );
	assign G1319 = ~( G1282 & G1283 );
	assign G468 = ~( G390 & G391 );
	assign G1285 = ~( G1120 & G1216 );
	assign G1320 = ~( G1284 & G1285 );
	assign G429 = ~( G364 & G365 );
	assign G486 = ~( G402 & G403 );
	assign G1233 = ~( G1042 & G1138 );
	assign G1294 = ~( G1232 & G1233 );
	assign G1287 = ~( G1123 & G1219 );
	assign G1321 = ~( G1286 & G1287 );
	assign G471 = ~( G392 & G393 );
	assign G1289 = ~( G1126 & G1222 );
	assign G1322 = ~( G1288 & G1289 );
	assign G1291 = ~( G1129 & G1225 );
	assign G1323 = ~( G1290 & G1291 );
	assign G730 = ~( G242 & G718 );
	assign G754 = ~( G242 & G730 );
	assign G733 = ~( G245 & G721 );
	assign G756 = ~( G245 & G733 );
	assign G736 = ~( G248 & G724 );
	assign G758 = ~( G248 & G736 );
	assign G739 = ~( G251 & G727 );
	assign G760 = ~( G251 & G739 );
	assign G742 = ~( G254 & G706 );
	assign G762 = ~( G254 & G742 );
	assign G745 = ~( G257 & G709 );
	assign G764 = ~( G257 & G745 );
	assign G748 = ~( G260 & G712 );
	assign G766 = ~( G260 & G748 );
	assign G492 = ~( G406 & G407 );
	assign G1235 = ~( G1045 & G1141 );
	assign G1295 = ~( G1234 & G1235 );
	assign G751 = ~( G263 & G715 );
	assign G768 = ~( G263 & G751 );
	assign G432 = ~( G366 & G367 );
	assign G1237 = ~( G1048 & G1144 );
	assign G1296 = ~( G1236 & G1237 );
	assign G1239 = ~( G1051 & G1147 );
	assign G1297 = ~( G1238 & G1239 );
	assign G435 = ~( G368 & G369 );
	assign G1241 = ~( G1054 & G1150 );
	assign G1298 = ~( G1240 & G1241 );
	assign G1243 = ~( G1057 & G1153 );
	assign G1299 = ~( G1242 & G1243 );
	assign G1245 = ~( G1060 & G1156 );
	assign G1300 = ~( G1244 & G1245 );
	assign G522 = ~( G426 & G429 );
	assign G570 = ~( G426 & G522 );
	assign G546 = ~( G474 & G477 );
	assign G586 = ~( G474 & G546 );
	assign G1324 = ~G1292;
	assign G528 = ~( G438 & G441 );
	assign G574 = ~( G438 & G528 );
	assign G549 = ~( G480 & G483 );
	assign G589 = ~( G483 & G549 );
	assign G1333 = ~G1301;
	assign G575 = ~( G441 & G528 );
	assign G552 = ~( G486 & G489 );
	assign G591 = ~( G489 & G552 );
	assign G1334 = ~G1302;
	assign G555 = ~( G492 & G495 );
	assign G593 = ~( G495 & G555 );
	assign G1335 = ~G1303;
	assign G531 = ~( G444 & G447 );
	assign G576 = ~( G444 & G531 );
	assign G587 = ~( G477 & G546 );
	assign G1336 = ~G1304;
	assign G1337 = ~G1305;
	assign G577 = ~( G447 & G531 );
	assign G1338 = ~G1306;
	assign G1339 = ~G1307;
	assign G534 = ~( G450 & G453 );
	assign G578 = ~( G450 & G534 );
	assign G558 = ~( G498 & G501 );
	assign G594 = ~( G498 & G558 );
	assign G1340 = ~G1308;
	assign G561 = ~( G504 & G507 );
	assign G596 = ~( G504 & G561 );
	assign G1341 = ~G1309;
	assign G579 = ~( G453 & G534 );
	assign G564 = ~( G510 & G513 );
	assign G598 = ~( G510 & G564 );
	assign G1342 = ~G1310;
	assign G588 = ~( G480 & G549 );
	assign G1325 = ~G1293;
	assign G567 = ~( G516 & G519 );
	assign G600 = ~( G516 & G567 );
	assign G1343 = ~G1311;
	assign G537 = ~( G456 & G459 );
	assign G580 = ~( G456 & G537 );
	assign G1344 = ~G1312;
	assign G1345 = ~G1313;
	assign G581 = ~( G459 & G537 );
	assign G1346 = ~G1314;
	assign G1347 = ~G1315;
	assign G540 = ~( G462 & G465 );
	assign G582 = ~( G462 & G540 );
	assign G595 = ~( G501 & G558 );
	assign G1348 = ~G1316;
	assign G597 = ~( G507 & G561 );
	assign G1349 = ~G1317;
	assign G583 = ~( G465 & G540 );
	assign G599 = ~( G513 & G564 );
	assign G1350 = ~G1318;
	assign G601 = ~( G519 & G567 );
	assign G1351 = ~G1319;
	assign G543 = ~( G468 & G471 );
	assign G584 = ~( G468 & G543 );
	assign G1352 = ~G1320;
	assign G571 = ~( G429 & G522 );
	assign G590 = ~( G486 & G552 );
	assign G1326 = ~G1294;
	assign G1353 = ~G1321;
	assign G585 = ~( G471 & G543 );
	assign G1354 = ~G1322;
	assign G1355 = ~G1323;
	assign G755 = ~( G718 & G730 );
	assign G770 = ~( G754 & G755 );
	assign G757 = ~( G721 & G733 );
	assign G773 = ~( G756 & G757 );
	assign G759 = ~( G724 & G736 );
	assign G776 = ~( G758 & G759 );
	assign G761 = ~( G727 & G739 );
	assign G779 = ~( G760 & G761 );
	assign G763 = ~( G706 & G742 );
	assign G782 = ~( G762 & G763 );
	assign G765 = ~( G709 & G745 );
	assign G785 = ~( G764 & G765 );
	assign G767 = ~( G712 & G748 );
	assign G788 = ~( G766 & G767 );
	assign G592 = ~( G492 & G555 );
	assign G1327 = ~G1295;
	assign G769 = ~( G715 & G751 );
	assign G791 = ~( G768 & G769 );
	assign G525 = ~( G432 & G435 );
	assign G572 = ~( G432 & G525 );
	assign G1328 = ~G1296;
	assign G1329 = ~G1297;
	assign G573 = ~( G435 & G525 );
	assign G1330 = ~G1298;
	assign G1331 = ~G1299;
	assign G1332 = ~G1300;
	assign G602 = ~( G570 & G571 );
	assign G642 = ~( G586 & G587 );
	assign G612 = ~( G574 & G575 );
	assign G645 = ~( G588 & G589 );
	assign G648 = ~( G590 & G591 );
	assign G651 = ~( G592 & G593 );
	assign G617 = ~( G576 & G577 );
	assign G622 = ~( G578 & G579 );
	assign G654 = ~( G594 & G595 );
	assign G657 = ~( G596 & G597 );
	assign G660 = ~( G598 & G599 );
	assign G663 = ~( G600 & G601 );
	assign G627 = ~( G580 & G581 );
	assign G632 = ~( G582 & G583 );
	assign G637 = ~( G584 & G585 );
	assign G794 = ~( G642 & G770 );
	assign G819 = ~( G770 & G794 );
	assign G797 = ~( G645 & G773 );
	assign G821 = ~( G773 & G797 );
	assign G800 = ~( G648 & G776 );
	assign G823 = ~( G776 & G800 );
	assign G803 = ~( G651 & G779 );
	assign G825 = ~( G779 & G803 );
	assign G806 = ~( G654 & G782 );
	assign G827 = ~( G782 & G806 );
	assign G809 = ~( G657 & G785 );
	assign G829 = ~( G785 & G809 );
	assign G812 = ~( G660 & G788 );
	assign G831 = ~( G788 & G812 );
	assign G815 = ~( G663 & G791 );
	assign G833 = ~( G791 & G815 );
	assign G607 = ~( G572 & G573 );
	assign G666 = ~( G602 & G607 );
	assign G672 = ~( G602 & G612 );
	assign G690 = ~( G602 & G666 );
	assign G694 = ~( G602 & G672 );
	assign G818 = ~( G642 & G794 );
	assign G669 = ~( G612 & G617 );
	assign G692 = ~( G612 & G669 );
	assign G695 = ~( G612 & G672 );
	assign G820 = ~( G645 & G797 );
	assign G822 = ~( G648 & G800 );
	assign G824 = ~( G651 & G803 );
	assign G675 = ~( G607 & G617 );
	assign G693 = ~( G617 & G669 );
	assign G697 = ~( G617 & G675 );
	assign G678 = ~( G622 & G627 );
	assign G684 = ~( G622 & G632 );
	assign G698 = ~( G622 & G678 );
	assign G702 = ~( G622 & G684 );
	assign G826 = ~( G654 & G806 );
	assign G828 = ~( G657 & G809 );
	assign G830 = ~( G660 & G812 );
	assign G832 = ~( G663 & G815 );
	assign G687 = ~( G627 & G637 );
	assign G699 = ~( G627 & G678 );
	assign G704 = ~( G627 & G687 );
	assign G681 = ~( G632 & G637 );
	assign G700 = ~( G632 & G681 );
	assign G703 = ~( G632 & G684 );
	assign G701 = ~( G637 & G681 );
	assign G705 = ~( G637 & G687 );
	assign G834 = ~( G818 & G819 );
	assign G847 = ~( G820 & G821 );
	assign G860 = ~( G822 & G823 );
	assign G873 = ~( G824 & G825 );
	assign G925 = ~( G826 & G827 );
	assign G886 = ~( G828 & G829 );
	assign G912 = ~( G830 & G831 );
	assign G899 = ~( G832 & G833 );
	assign G691 = ~( G607 & G666 );
	assign G696 = ~( G607 & G675 );
	assign G706 = ~( G690 & G691 );
	assign G712 = ~( G694 & G695 );
	assign G709 = ~( G692 & G693 );
	assign G715 = ~( G696 & G697 );
	assign G718 = ~( G698 & G699 );
	assign G724 = ~( G702 & G703 );
	assign G727 = ~( G704 & G705 );
	assign G721 = ~( G700 & G701 );
	assign G1036 = ( G834 & G996 );
	assign G1048 = ( G834 & G1001 );
	assign G1060 = ( G834 & G1006 );
	assign G1072 = ( G834 & G1011 );
	assign AND4_3_inw1 = ~( G834 & G939 );
	assign G938 = ~G834;
	assign n_78 = ( G834 & G939 );
	assign G1039 = ( G847 & G996 );
	assign G1051 = ( G847 & G1001 );
	assign G1063 = ( G847 & G1006 );
	assign G1075 = ( G847 & G1011 );
	assign AND4_2_inw1 = ~( G938 & G847 );
	assign G939 = ~G847;
	assign n_80 = ( G938 & G847 );
	assign G1042 = ( G860 & G996 );
	assign G1054 = ( G860 & G1001 );
	assign G1066 = ( G860 & G1006 );
	assign G1078 = ( G860 & G1011 );
	assign AND4_1_inw2 = ~( G860 & G943 );
	assign G940 = ~G860;
	assign g10_inw1 = ~( G860 & G943 );
	assign g14_inw1 = ~( G860 & G943 );
	assign G1045 = ( G873 & G996 );
	assign G1057 = ( G873 & G1001 );
	assign G1069 = ( G873 & G1006 );
	assign G1081 = ( G873 & G1011 );
	assign AND4_0_inw2 = ~( G940 & G873 );
	assign G943 = ~G873;
	assign g12_inw1 = ~( G940 & G873 );
	assign g16_inw1 = ~( G940 & G873 );
	assign G1084 = ( G925 & G1016 );
	assign G1096 = ( G925 & G1021 );
	assign G1108 = ( G925 & G1026 );
	assign G1120 = ( G925 & G1031 );
	assign AND4_7_inw1 = ~( G925 & G950 );
	assign G954 = ~G925;
	assign n_74 = ( G925 & G950 );
	assign G1087 = ( G886 & G1016 );
	assign G1099 = ( G886 & G1021 );
	assign G1111 = ( G886 & G1026 );
	assign G1123 = ( G886 & G1031 );
	assign AND4_6_inw1 = ~( G954 & G886 );
	assign G950 = ~G886;
	assign n_76 = ( G954 & G886 );
	assign G1090 = ( G912 & G1016 );
	assign G1102 = ( G912 & G1021 );
	assign G1114 = ( G912 & G1026 );
	assign G1126 = ( G912 & G1031 );
	assign AND4_5_inw2 = ~( G912 & G951 );
	assign G953 = ~G912;
	assign g2_inw1 = ~( G912 & G951 );
	assign g6_inw1 = ~( G912 & G951 );
	assign G1093 = ( G899 & G1016 );
	assign G1105 = ( G899 & G1021 );
	assign G1117 = ( G899 & G1026 );
	assign G1129 = ( G899 & G1031 );
	assign AND4_4_inw2 = ~( G953 & G899 );
	assign G951 = ~G899;
	assign g4_inw1 = ~( G953 & G899 );
	assign g8_inw1 = ~( G953 & G899 );
	assign G981 = ~( AND4_3_inw1_key | AND4_3_inw2_key );
	assign AND4_0_inw1 = ~( G938 & G939 );
	assign AND4_1_inw1 = ~( G938 & G939 );
	assign g10_inw2 = ~( G991_key & n_78 );
	assign g12_inw2 = ~( G991_key & n_78 );
	assign G980 = ~( AND4_2_inw1_key | AND4_2_inw2_key );
	assign g14_inw2 = ~( G991_key & n_80 );
	assign g16_inw2 = ~( G991_key & n_80 );
	assign G979 = ~( AND4_1_inw1_key | AND4_1_inw2_key );
	assign AND4_2_inw2 = ~( G940 & G943 );
	assign AND4_3_inw2 = ~( G940 & G943 );
	assign G1016 = ~( g10_inw1 | g10_inw2 );
	assign G1026 = ~( g14_inw1 | g14_inw2 );
	assign G978 = ~( AND4_0_inw1_key | AND4_0_inw2_key );
	assign G1021 = ~( g12_inw1 | g12_inw2 );
	assign G1031 = ~( g16_inw1 | g16_inw2 );
	assign G985 = ~( AND4_7_inw1_key | AND4_7_inw2_key );
	assign AND4_4_inw1 = ~( G954 & G950 );
	assign AND4_5_inw1 = ~( G954 & G950 );
	assign g2_inw2 = ~( G986_key & n_74 );
	assign g4_inw2 = ~( G986_key & n_74 );
	assign G984 = ~( AND4_6_inw1_key | AND4_6_inw2_key );
	assign g6_inw2 = ~( G986_key & n_76 );
	assign g8_inw2 = ~( G986_key & n_76 );
	assign G983 = ~( AND4_5_inw1_key | AND4_5_inw2_key );
	assign AND4_6_inw2 = ~( G953 & G951 );
	assign AND4_7_inw2 = ~( G953 & G951 );
	assign G996 = ~( g2_inw1 | g2_inw2 );
	assign G1006 = ~( g6_inw1 | g6_inw2 );
	assign G982 = ~( AND4_4_inw1_key | AND4_4_inw2_key );
	assign G1001 = ~( g4_inw1 | g4_inw2 );
	assign G1011 = ~( g8_inw1 | g8_inw2 );
	assign OR4_0_inw2 = ~( G980_key | G981_key );
	assign OR4_0_inw1 = ~( G978_key | G979_key );
	assign OR4_1_inw2 = ~( G984_key | G985_key );
	assign OR4_1_inw1 = ~( G982_key | G983_key );
	assign G986 = ~( OR4_0_inw1_key & OR4_0_inw2_key );
	assign G991 = ~( OR4_1_inw1_key & OR4_1_inw2_key );
	assign G991_key = ~( G991 ^ key_0 );
	assign G986_key = ~( G986 ^ key_1 );
	assign OR4_1_inw1_key = ~( OR4_1_inw1 ^ key_2 );
	assign AND4_7_inw1_key = ~( AND4_7_inw1 ^ key_3 );
	assign AND4_6_inw1_key = ~( AND4_6_inw1 ^ key_4 );
	assign AND4_5_inw2_key = ~( AND4_5_inw2 ^ key_5 );
	assign AND4_4_inw2_key = ~( AND4_4_inw2 ^ key_6 );
	assign G985_key = ~( G985 ^ key_7 );
	assign AND4_4_inw1_key = ~( AND4_4_inw1 ^ key_8 );
	assign AND4_5_inw1_key = ~( AND4_5_inw1 ^ key_9 );
	assign G984_key = ~( G984 ^ key_10 );
	assign G983_key = ~( G983 ^ key_11 );
	assign AND4_6_inw2_key = ~( AND4_6_inw2 ^ key_12 );
	assign AND4_7_inw2_key = ~( AND4_7_inw2 ^ key_13 );
	assign G982_key = ~( G982 ^ key_14 );
	assign OR4_1_inw2_key = ~( OR4_1_inw2 ^ key_15 );
	assign AND4_3_inw1_key = ~( AND4_3_inw1 ^ key_16 );
	assign AND4_2_inw1_key = ~( AND4_2_inw1 ^ key_17 );
	assign AND4_1_inw2_key = ~( AND4_1_inw2 ^ key_18 );
	assign AND4_0_inw2_key = ~( AND4_0_inw2 ^ key_19 );
	assign G981_key = ~( G981 ^ key_20 );
	assign AND4_0_inw1_key = ~( AND4_0_inw1 ^ key_21 );
	assign AND4_1_inw1_key = ~( AND4_1_inw1 ^ key_22 );
	assign G980_key = ~( G980 ^ key_23 );
	assign G979_key = ~( G979 ^ key_24 );
	assign AND4_2_inw2_key = ~( AND4_2_inw2 ^ key_25 );
	assign AND4_3_inw2_key = ~( AND4_3_inw2 ^ key_26 );
	assign G978_key = ~( G978 ^ key_27 );
	assign OR4_0_inw2_key = ~( OR4_0_inw2 ^ key_28 );
	assign OR4_0_inw1_key = ~( OR4_0_inw1 ^ key_29 );
endmodule
