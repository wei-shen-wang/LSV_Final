module c880(N1, N101, N106, N111, N116, N121, N126, N13, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N17, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N26, N260, N261, N267, N268, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N8, N80, N85, N86, N87, N88, N89, N90, N91, N96, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880);
	input N1, N101, N106, N111, N116, N121, N126, N13, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N17, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N26, N260, N261, N267, N268, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N8, N80, N85, N86, N87, N88, N89, N90, N91, N96;
	output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
	wire N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, AND3_4_inw1, N483, NAND4_1_inw1, NAND4_2_inw1, NAND4_5_inw1, NAND4_6_inw1, N309, NAND4_1_inw2, NAND4_2_inw2, NAND4_6_inw2, N317, N323, NAND3_117_invw, NAND4_5_inw2, N322, g13_inw2, AND3_3_inw1, AND3_10_inw1, AND3_11_inw1, AND3_12_inw1, N285, AND3_16_inw1, AND3_17_inw1, N390, N388, N294, N296, n_92, N316, N447, N427, n_95, AND3_14_inw1, AND3_15_inw1, N319, NAND4_116_inw1, n_87, n_91, n_88, g8_inw1, n_89, N287, N389, N293, N295, N391, N298, N355, N423, N332, N502, N301, N302, N333, N504, N334, N506, N303, N304, N335, N508, N336, N511, N305, N306, N338, N513, N340, N515, N307, N308, N517, N498, N518, N499, N519, N500, N501, N318, N475, N510, N477, N512, N479, N514, N481, N516, NAND4_116_inw2, N522, N324, N590, N325, N593, N523, N597, N600, N524, N326, N606, N327, N609, N525, N616, N619, N526, N328, N625, N329, N628, N527, N632, N635, N330, N528, N641, N331, N644, N529, N651, N654, N520, N521, N417, N794, N808, N809, N810, N836, N851, N852, N853, N736, N739, N742, N745, N748, N751, N754, N759, N737, N740, N743, N746, N749, N752, N755, N760, N596, N605, N615, N624, N631, N640, N650, N659, N337, N339, N341, N758, N732, NAND3_255_invw, NAND4_256_inw2, N757, g9_inw2, n_96, NAND4_1_invw, NAND4_2_invw, NAND4_5_invw, NAND4_6_invw, N536, N538, N375, N443, N476, N349, N343, N419, N352, N422, g8_inw2, N537, AND3_113_inw1, NAND3_117_inw1, n_93, g13_inw1, NAND4_116_invw, g1_inw1, N400, g1_inw2, n_94, N420, N421, N450, N860, N357, N861, N845, N360, N826, N539, N827, N540, N363, N828, N541, N805, N542, N366, N543, N530, N544, N533, N503, N505, N507, N509, N669, N376, N665, N849, N662, N841, N677, N673, NAND4_325_inw1, N670, N765, NAND3_288_inw1, NAND4_324_inw1, N686, N379, N682, NAND3_326_inw1, N678, N764, NAND3_323_inw1, N696, N692, N822, N687, N812, NAND4_324_inw2, N704, N382, N700, N796, N697, N795, NAND4_341_inw2, N708, NAND4_295_inw1, N705, N762, NAND3_285_inw1, NAND4_256_inw1, N385, NAND4_342_inw2, N717, NAND3_297_inw1, N713, N761, NAND3_255_inw1, NAND4_321_inw2, N727, N782, N722, N547, N859, N769, N770, N771, N772, N777, N781, N785, N787, N712, N721, N731, N786, N733, NAND4_256_invw, N488, N269, N270, N279, N280, N553, N561, N448, N446, N410, N557, g9_inw1, N442, N350, NAND3_371_inw1, N406, N404, NAND3_372_inw1, NAND3_357_inw1, N405, NAND3_340_inw1, N565, NAND4_341_inw1, N569, N409, N407, NAND4_342_inw1, N573, NAND4_321_inw1, N577, N408, N581, N552, N550, N587, N585, N551, NAND3_370_invw, N413, N411, N831, N830, N866, NAND3_371_invw, N833, N832, NAND4_325_invw, NAND3_288_invw, NAND4_324_invw, NAND3_372_invw, N412, N835, N834, NAND3_326_invw, NAND3_323_invw, NAND3_357_invw, N807, N806, NAND3_340_invw, N416, N414, N789, N788, NAND4_341_invw, N791, N790, NAND4_295_invw, NAND3_285_invw, N415, NAND4_342_invw, N793, N792, NAND3_297_invw, NAND4_321_invw, N586, NAND3_370_inw1, N734, N418, N347, n_90, N466, N449, N460, N425, N463, N426, N767, N588, N768, N589, N878, N492, N444, N842, N879, N843, N815, N766, N814, N880, N844, N819, N813, N874, N825, N863, N495, N445, N802, N864, N803, N773, N763, N865, N804, N778, N850, NAND4_295_inw2, NAND4_325_inw2;
	assign AND3_4_inw1 = ~( N1 & N26 );
	assign N483 = ~( N443 & N1 );
	assign NAND4_1_inw1 = ~( N1 & N8 );
	assign NAND4_2_inw1 = ~( N1 & N26 );
	assign NAND4_5_inw1 = ~( N1 & N8 );
	assign NAND4_6_inw1 = ~( N1 & N8 );
	assign N309 = ( N8 & N138 );
	assign NAND4_1_inw2 = ~( N13 & N17 );
	assign NAND4_2_inw2 = ~( N13 & N17 );
	assign NAND4_6_inw2 = ~( N13 & N55 );
	assign N317 = ( N17 & N138 );
	assign N323 = ( N17 & N42 );
	assign NAND3_117_invw = ~( NAND3_117_inw1 | N17 );
	assign NAND4_5_inw2 = ~( N51 & N17 );
	assign N322 = ~( N17 | N42 );
	assign g13_inw2 = ~( N17 & N287 );
	assign AND3_3_inw1 = ~( N29 & N36 );
	assign AND3_10_inw1 = ~( N29 & N75 );
	assign AND3_11_inw1 = ~( N29 & N75 );
	assign AND3_12_inw1 = ~( N29 & N36 );
	assign N285 = ~( N29 & N68 );
	assign AND3_16_inw1 = ~( N59 & N36 );
	assign AND3_17_inw1 = ~( N59 & N36 );
	assign N390 = ~( AND3_3_inw1 | N42 );
	assign N388 = ~( AND3_11_inw1 | N42 );
	assign N294 = ~( AND3_15_inw1 | N42 );
	assign N296 = ~( AND3_17_inw1 | N42 );
	assign n_92 = ( N42 & N68 );
	assign N316 = ( N51 & N138 );
	assign N447 = ~( AND3_4_inw1 | N51 );
	assign N427 = ~( AND3_113_inw1 | N55 );
	assign n_95 = ~N55;
	assign AND3_14_inw1 = ~( N59 & N75 );
	assign AND3_15_inw1 = ~( N59 & N75 );
	assign N319 = ~( N59 & N156 );
	assign NAND4_116_inw1 = ~( N375 & N59 );
	assign n_87 = ~N59;
	assign n_91 = ( n_90 & N59 );
	assign n_88 = ~N68;
	assign g8_inw1 = ~( N72 & N73 );
	assign n_89 = ~N74;
	assign N287 = ~( AND3_10_inw1 | N80 );
	assign N389 = ~( AND3_12_inw1 | N80 );
	assign N293 = ~( AND3_14_inw1 | N80 );
	assign N295 = ~( AND3_16_inw1 | N80 );
	assign N391 = ( N85 & N86 );
	assign N298 = ( N87 | N88 );
	assign N355 = ~( N89 & N298 );
	assign N423 = ( N90 & N298 );
	assign N332 = ( N210 & N91 );
	assign N502 = ( N91 & N466 );
	assign N301 = ~( N91 & N96 );
	assign N302 = ( N91 | N96 );
	assign N333 = ( N210 & N96 );
	assign N504 = ( N96 & N466 );
	assign N334 = ( N210 & N101 );
	assign N506 = ( N101 & N466 );
	assign N303 = ~( N101 & N106 );
	assign N304 = ( N101 | N106 );
	assign N335 = ( N210 & N106 );
	assign N508 = ( N106 & N466 );
	assign N336 = ( N210 & N111 );
	assign N511 = ( N111 & N466 );
	assign N305 = ~( N111 & N116 );
	assign N306 = ( N111 | N116 );
	assign N338 = ( N210 & N116 );
	assign N513 = ( N116 & N466 );
	assign N340 = ( N210 & N121 );
	assign N515 = ( N121 & N466 );
	assign N307 = ~( N121 & N126 );
	assign N308 = ( N121 | N126 );
	assign N517 = ( N126 & N466 );
	assign N498 = ~( N130 & N460 );
	assign N518 = ~( N130 & N492 );
	assign N499 = ( N130 | N460 );
	assign N519 = ( N130 | N492 );
	assign N500 = ~( N463 & N135 );
	assign N501 = ( N463 | N135 );
	assign N318 = ( N152 & N138 );
	assign N475 = ( N143 & N427 );
	assign N510 = ( N143 & N483 );
	assign N477 = ( N146 & N427 );
	assign N512 = ( N146 & N483 );
	assign N479 = ( N149 & N427 );
	assign N514 = ( N149 & N483 );
	assign N481 = ( N153 & N427 );
	assign N516 = ( N153 & N483 );
	assign NAND4_116_inw2 = ~( N156 & N447 );
	assign N522 = ( N400 & N159 );
	assign N324 = ~( N159 & N165 );
	assign N590 = ~( N553 & N159 );
	assign N325 = ( N159 | N165 );
	assign N593 = ( N553 | N159 );
	assign N523 = ( N400 & N165 );
	assign N597 = ~( N557 & N165 );
	assign N600 = ( N557 | N165 );
	assign N524 = ( N400 & N171 );
	assign N326 = ~( N171 & N177 );
	assign N606 = ~( N561 & N171 );
	assign N327 = ( N171 | N177 );
	assign N609 = ( N561 | N171 );
	assign N525 = ( N400 & N177 );
	assign N616 = ~( N565 & N177 );
	assign N619 = ( N565 | N177 );
	assign N526 = ( N400 & N183 );
	assign N328 = ~( N183 & N189 );
	assign N625 = ~( N569 & N183 );
	assign N329 = ( N183 | N189 );
	assign N628 = ( N569 | N183 );
	assign N527 = ~( N400 & N189 );
	assign N632 = ~( N573 & N189 );
	assign N635 = ( N573 | N189 );
	assign N330 = ~( N195 & N201 );
	assign N528 = ~( N400 & N195 );
	assign N641 = ~( N577 & N195 );
	assign N331 = ( N195 | N201 );
	assign N644 = ( N577 | N195 );
	assign N529 = ~( N400 & N201 );
	assign N651 = ~( N581 & N201 );
	assign N654 = ( N581 | N201 );
	assign N520 = ~( N495 & N207 );
	assign N521 = ( N495 | N207 );
	assign N417 = ( N210 & N268 );
	assign N794 = ( N219 & N786 );
	assign N808 = ( N219 & N802 );
	assign N809 = ( N219 & N803 );
	assign N810 = ( N219 & N804 );
	assign N836 = ( N219 & N825 );
	assign N851 = ( N219 & N842 );
	assign N852 = ( N219 & N843 );
	assign N853 = ( N219 & N844 );
	assign N736 = ( N228 & N665 );
	assign N739 = ( N228 & N673 );
	assign N742 = ( N228 & N682 );
	assign N745 = ( N228 & N692 );
	assign N748 = ( N228 & N700 );
	assign N751 = ( N228 & N708 );
	assign N754 = ( N228 & N717 );
	assign N759 = ( N228 & N727 );
	assign N737 = ( N237 & N662 );
	assign N740 = ( N237 & N670 );
	assign N743 = ( N237 & N678 );
	assign N746 = ( N237 & N687 );
	assign N749 = ( N237 & N697 );
	assign N752 = ( N237 & N705 );
	assign N755 = ( N237 & N713 );
	assign N760 = ( N237 & N722 );
	assign N596 = ( N246 & N553 );
	assign N605 = ( N246 & N557 );
	assign N615 = ( N246 & N561 );
	assign N624 = ( N246 & N565 );
	assign N631 = ( N246 & N569 );
	assign N640 = ( N246 & N573 );
	assign N650 = ( N246 & N577 );
	assign N659 = ( N246 & N581 );
	assign N337 = ( N255 & N259 );
	assign N339 = ( N255 & N260 );
	assign N341 = ( N255 & N267 );
	assign N758 = ( N727 & N261 );
	assign N732 = ~( N654 & N261 );
	assign NAND3_255_invw = ~( NAND3_255_inw1 | N261 );
	assign NAND4_256_inw2 = ~( N654 & N261 );
	assign N757 = ~( N727 | N261 );
	assign g9_inw2 = ~( n_95 | N268 );
	assign n_96 = ~N268;
	assign NAND4_1_invw = ~( NAND4_1_inw1 | NAND4_1_inw2 );
	assign NAND4_2_invw = ~( NAND4_2_inw1 | NAND4_2_inw2 );
	assign NAND4_5_invw = ~( NAND4_5_inw1 | NAND4_5_inw2 );
	assign NAND4_6_invw = ~( NAND4_6_inw1 | NAND4_6_inw2 );
	assign N536 = ~( N309 | N502 );
	assign N538 = ~( N317 | N506 );
	assign N375 = ~( N322 | N323 );
	assign N443 = ~NAND3_117_invw;
	assign N476 = ~( g13_inw1 | g13_inw2 );
	assign N349 = ( N280 | N285 );
	assign N343 = ~N390;
	assign N419 = ( N270 | N390 );
	assign N352 = ~N294;
	assign N422 = ~N296;
	assign g8_inw2 = ~( n_91 & n_92 );
	assign N537 = ~( N316 | N504 );
	assign AND3_113_inw1 = ~( N319 & N447 );
	assign NAND3_117_inw1 = ~( N447 & N319 );
	assign n_93 = ~N447;
	assign g13_inw1 = ~( n_96 & N447 );
	assign NAND4_116_invw = ~( NAND4_116_inw1 | NAND4_116_inw2 );
	assign g1_inw1 = ~( n_87 | n_88 );
	assign N400 = ~( g8_inw1 | g8_inw2 );
	assign g1_inw2 = ~( n_89 | N280 );
	assign n_94 = ~N287;
	assign N420 = ~N293;
	assign N421 = ~N295;
	assign N450 = ~N355;
	assign N860 = ~( N332 | N852 );
	assign N357 = ~( N301 & N302 );
	assign N861 = ~( N333 | N853 );
	assign N845 = ~( N334 | N836 );
	assign N360 = ~( N303 & N304 );
	assign N826 = ~( N335 | N808 );
	assign N539 = ~( N318 | N508 );
	assign N827 = ~( N336 | N809 );
	assign N540 = ~( N510 | N511 );
	assign N363 = ~( N305 & N306 );
	assign N828 = ~( N338 | N810 );
	assign N541 = ~( N512 | N513 );
	assign N805 = ~( N340 | N794 );
	assign N542 = ~( N514 | N515 );
	assign N366 = ~( N307 & N308 );
	assign N543 = ~( N516 | N517 );
	assign N530 = ~( N498 & N499 );
	assign N544 = ~( N518 & N519 );
	assign N533 = ~( N500 & N501 );
	assign N503 = ~( N475 | N476 );
	assign N505 = ~( N477 | N476 );
	assign N507 = ~( N479 | N476 );
	assign N509 = ~( N481 | N476 );
	assign N669 = ~( N596 | N522 );
	assign N376 = ~( N324 & N325 );
	assign N665 = ( N593 & N590 );
	assign N849 = ( N590 & N841 );
	assign N662 = ~N590;
	assign N841 = ~( N815 & N593 );
	assign N677 = ~( N605 | N523 );
	assign N673 = ( N600 & N597 );
	assign NAND4_325_inw1 = ~( N597 & N765 );
	assign N670 = ~N597;
	assign N765 = ~( N600 & N678 );
	assign NAND3_288_inw1 = ~( N600 & N609 );
	assign NAND4_324_inw1 = ~( N600 & N609 );
	assign N686 = ~( N615 | N524 );
	assign N379 = ~( N326 & N327 );
	assign N682 = ( N609 & N606 );
	assign NAND3_326_inw1 = ~( N606 & N764 );
	assign N678 = ~N606;
	assign N764 = ~( N609 & N687 );
	assign NAND3_323_inw1 = ~( N609 & N619 );
	assign N696 = ~( N624 | N525 );
	assign N692 = ( N619 & N616 );
	assign N822 = ~( N616 & N812 );
	assign N687 = ~N616;
	assign N812 = ~( N619 & N796 );
	assign NAND4_324_inw2 = ~( N619 & N796 );
	assign N704 = ~( N631 | N526 );
	assign N382 = ~( N328 & N329 );
	assign N700 = ( N628 & N625 );
	assign N796 = ~( N795 & N625 );
	assign N697 = ~N625;
	assign N795 = ~( N628 & N773 );
	assign NAND4_341_inw2 = ~( N712 & N527 );
	assign N708 = ( N635 & N632 );
	assign NAND4_295_inw1 = ~( N632 & N762 );
	assign N705 = ~N632;
	assign N762 = ~( N635 & N713 );
	assign NAND3_285_inw1 = ~( N635 & N644 );
	assign NAND4_256_inw1 = ~( N635 & N644 );
	assign N385 = ~( N330 & N331 );
	assign NAND4_342_inw2 = ~( N721 & N528 );
	assign N717 = ( N644 & N641 );
	assign NAND3_297_inw1 = ~( N641 & N761 );
	assign N713 = ~N641;
	assign N761 = ~( N644 & N722 );
	assign NAND3_255_inw1 = ~( N644 & N654 );
	assign NAND4_321_inw2 = ~( N731 & N529 );
	assign N727 = ( N654 & N651 );
	assign N782 = ~( N651 & N732 );
	assign N722 = ~N651;
	assign N547 = ~( N520 & N521 );
	assign N859 = ~( N417 | N851 );
	assign N769 = ~( N736 | N737 );
	assign N770 = ~( N739 | N740 );
	assign N771 = ~( N742 | N743 );
	assign N772 = ~( N745 | N746 );
	assign N777 = ~( N748 | N749 );
	assign N781 = ~( N751 | N752 );
	assign N785 = ~( N754 | N755 );
	assign N787 = ~( N759 | N760 );
	assign N712 = ~( N337 | N640 );
	assign N721 = ~( N339 | N650 );
	assign N731 = ~( N341 | N659 );
	assign N786 = ~( N757 | N758 );
	assign N733 = ~NAND3_255_invw;
	assign NAND4_256_invw = ~( NAND4_256_inw1 | NAND4_256_inw2 );
	assign N488 = ~( g9_inw1 & g9_inw2 );
	assign N269 = ~NAND4_1_invw;
	assign N270 = ~NAND4_2_invw;
	assign N279 = ~NAND4_5_invw;
	assign N280 = ~NAND4_6_invw;
	assign N553 = ~( N536 & N503 );
	assign N561 = ~( N538 & N507 );
	assign N448 = ~N349;
	assign N446 = ( N270 | N343 );
	assign N410 = ~( N347 & N352 );
	assign N557 = ~( N537 & N505 );
	assign g9_inw1 = ~( n_93 | n_94 );
	assign N442 = ~NAND4_116_invw;
	assign N350 = ~( g1_inw1 & g1_inw2 );
	assign NAND3_371_inw1 = ~( N860 & N770 );
	assign N406 = ( N357 & N360 );
	assign N404 = ~N357;
	assign NAND3_372_inw1 = ~( N861 & N771 );
	assign NAND3_357_inw1 = ~( N845 & N772 );
	assign N405 = ~N360;
	assign NAND3_340_inw1 = ~( N826 & N777 );
	assign N565 = ~( N539 & N509 );
	assign NAND4_341_inw1 = ~( N827 & N781 );
	assign N569 = ~( N488 & N540 );
	assign N409 = ( N363 & N366 );
	assign N407 = ~N363;
	assign NAND4_342_inw1 = ~( N828 & N785 );
	assign N573 = ~( N488 & N541 );
	assign NAND4_321_inw1 = ~( N805 & N787 );
	assign N577 = ~( N488 & N542 );
	assign N408 = ~N366;
	assign N581 = ~( N488 & N543 );
	assign N552 = ( N530 & N533 );
	assign N550 = ~N530;
	assign N587 = ( N544 & N547 );
	assign N585 = ~N544;
	assign N551 = ~N533;
	assign NAND3_370_invw = ~( NAND3_370_inw1 | N669 );
	assign N413 = ( N376 & N379 );
	assign N411 = ~N376;
	assign N831 = ( N665 & N815 );
	assign N830 = ~( N665 | N815 );
	assign N866 = ~N849;
	assign NAND3_371_invw = ~( NAND3_371_inw1 | N677 );
	assign N833 = ( N673 & N819 );
	assign N832 = ~( N673 | N819 );
	assign NAND4_325_invw = ~( NAND4_325_inw1 | NAND4_325_inw2 );
	assign NAND3_288_invw = ~( NAND3_288_inw1 | N687 );
	assign NAND4_324_invw = ~( NAND4_324_inw1 | NAND4_324_inw2 );
	assign NAND3_372_invw = ~( NAND3_372_inw1 | N686 );
	assign N412 = ~N379;
	assign N835 = ( N682 & N822 );
	assign N834 = ~( N682 | N822 );
	assign NAND3_326_invw = ~( NAND3_326_inw1 | N813 );
	assign NAND3_323_invw = ~( NAND3_323_inw1 | N796 );
	assign NAND3_357_invw = ~( NAND3_357_inw1 | N696 );
	assign N807 = ( N692 & N796 );
	assign N806 = ~( N692 | N796 );
	assign NAND3_340_invw = ~( NAND3_340_inw1 | N704 );
	assign N416 = ( N382 & N385 );
	assign N414 = ~N382;
	assign N789 = ( N700 & N773 );
	assign N788 = ~( N700 | N773 );
	assign NAND4_341_invw = ~( NAND4_341_inw1 | NAND4_341_inw2 );
	assign N791 = ( N708 & N778 );
	assign N790 = ~( N708 | N778 );
	assign NAND4_295_invw = ~( NAND4_295_inw1 | NAND4_295_inw2 );
	assign NAND3_285_invw = ~( NAND3_285_inw1 | N722 );
	assign N415 = ~N385;
	assign NAND4_342_invw = ~( NAND4_342_inw1 | NAND4_342_inw2 );
	assign N793 = ( N717 & N782 );
	assign N792 = ~( N717 | N782 );
	assign NAND3_297_invw = ~( NAND3_297_inw1 | N733 );
	assign NAND4_321_invw = ~( NAND4_321_inw1 | NAND4_321_inw2 );
	assign N586 = ~N547;
	assign NAND3_370_inw1 = ~( N859 & N769 );
	assign N734 = ~NAND4_256_invw;
	assign N418 = ~N269;
	assign N347 = ~N279;
	assign n_90 = ~N280;
	assign N466 = ~( N442 & N410 );
	assign N449 = ~N350;
	assign N460 = ~( N406 | N425 );
	assign N425 = ( N404 & N405 );
	assign N463 = ~( N409 | N426 );
	assign N426 = ( N407 & N408 );
	assign N767 = ~( N552 | N588 );
	assign N588 = ( N550 & N551 );
	assign N768 = ~( N587 | N589 );
	assign N589 = ( N585 & N586 );
	assign N878 = ~NAND3_370_invw;
	assign N492 = ~( N413 | N444 );
	assign N444 = ( N411 & N412 );
	assign N842 = ~( N830 | N831 );
	assign N879 = ~NAND3_371_invw;
	assign N843 = ~( N832 | N833 );
	assign N815 = ~NAND4_325_invw;
	assign N766 = ~NAND3_288_invw;
	assign N814 = ~NAND4_324_invw;
	assign N880 = ~NAND3_372_invw;
	assign N844 = ~( N834 | N835 );
	assign N819 = ~NAND3_326_invw;
	assign N813 = ~NAND3_323_invw;
	assign N874 = ~NAND3_357_invw;
	assign N825 = ~( N806 | N807 );
	assign N863 = ~NAND3_340_invw;
	assign N495 = ~( N416 | N445 );
	assign N445 = ( N414 & N415 );
	assign N802 = ~( N788 | N789 );
	assign N864 = ~NAND4_341_invw;
	assign N803 = ~( N790 | N791 );
	assign N773 = ~NAND4_295_invw;
	assign N763 = ~NAND3_285_invw;
	assign N865 = ~NAND4_342_invw;
	assign N804 = ~( N792 | N793 );
	assign N778 = ~NAND3_297_invw;
	assign N850 = ~NAND4_321_invw;
	assign NAND4_295_inw2 = ~( N763 & N734 );
	assign NAND4_325_inw2 = ~( N766 & N814 );
endmodule
