module c6288(N1, N103, N120, N137, N154, N171, N18, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N35, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N52, N528, N69, N86, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N545, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288);
	input N1, N103, N120, N137, N154, N171, N18, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N35, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N52, N528, N69, N86;
	output N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N545, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288;
	wire N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N546, N549, N552, N555, N558, N561, N564, N567, N570, N573, N576, N579, N582, N585, N588, N591, N594, N597, N600, N603, N606, N609, N612, N615, N618, N621, N624, N627, N630, N633, N636, N639, N642, N645, N648, N651, N654, N657, N660, N663, N666, N669, N672, N675, N678, N681, N684, N687, N690, N693, N696, N699, N702, N705, N708, N711, N714, N717, N720, N723, N726, N729, N732, N735, N738, N741, N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774, N777, N780, N783, N786, N789, N792, N795, N798, N801, N804, N807, N810, N813, N816, N819, N822, N825, N828, N831, N834, N837, N840, N843, N846, N849, N852, N855, N858, N861, N864, N867, N870, N873, N876, N879, N882, N885, N888, N891, N894, N897, N900, N903, N906, N909, N912, N915, N918, N921, N924, N927, N930, N933, N936, N939, N942, N945, N948, N951, N954, N957, N960, N963, N966, N969, N972, N975, N978, N981, N984, N987, N990, N993, N996, N999, N1002, N1005, N1008, N1011, N1014, N1017, N1020, N1023, N1026, N1029, N1032, N1035, N1038, N1041, N1044, N1047, N1050, N1053, N1056, N1059, N1062, N1065, N1068, N1071, N1074, N1077, N1080, N1083, N1086, N1089, N1092, N1095, N1098, N1101, N1104, N1107, N1110, N1113, N1116, N1119, N1122, N1125, N1128, N1131, N1134, N1137, N1140, N1143, N1146, N1149, N1152, N1155, N1158, N1161, N1164, N1167, N1170, N1173, N1176, N1179, N1182, N1185, N1188, N1191, N1194, N1197, N1200, N1203, N1206, N1209, N1212, N1215, N1218, N1221, N1224, N1227, N1230, N1233, N1236, N1239, N1242, N1245, N1248, N1251, N1254, N1257, N1260, N1263, N1266, N1269, N1272, N1275, N1278, N1281, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305, N1308, N1446, N1507, N1763, N1825, N2085, N2150, N2414, N2477, N2745, N2807, N3079, N3141, N3417, N3480, N3760, N3826, N4110, N4174, N4462, N4525, N4817, N4880, N5176, N5240, N5540, N5607, N5882, N5929, N6085, N6107, N1311, N1450, N1512, N1767, N1830, N2089, N2155, N2418, N2482, N2749, N2812, N3083, N3146, N3421, N3485, N3764, N3831, N4114, N4179, N4466, N4530, N4821, N4885, N5180, N5245, N5544, N5612, N5886, N5934, N6064, N6090, N1315, N1454, N1517, N1771, N1835, N2093, N2160, N2422, N2487, N2753, N2817, N3087, N3151, N3425, N3490, N3768, N3836, N4118, N4184, N4470, N4535, N4825, N4890, N5184, N5250, N5548, N5617, N5840, N5891, N6040, N6069, N1319, N1458, N1522, N1775, N1840, N2097, N2165, N2426, N2492, N2757, N2822, N3091, N3156, N3429, N3495, N3772, N3841, N4122, N4189, N4474, N4540, N4829, N4895, N5188, N5255, N5489, N5553, N5792, N5845, N6014, N6045, N1323, N1462, N1527, N1779, N1845, N2101, N2170, N2430, N2497, N2761, N2827, N3095, N3161, N3433, N3500, N3776, N3846, N4126, N4194, N4478, N4545, N4833, N4900, N5130, N5193, N5434, N5494, N5743, N5797, N5984, N6019, N1327, N1466, N1532, N1783, N1850, N2105, N2175, N2434, N2502, N2765, N2832, N3099, N3166, N3437, N3505, N3780, N3851, N4130, N4199, N4482, N4550, N4775, N4838, N5076, N5135, N5383, N5439, N5688, N5748, N5950, N5989, N1331, N1470, N1537, N1787, N1855, N2109, N2180, N2438, N2507, N2769, N2837, N3103, N3171, N3441, N3510, N3784, N3856, N4134, N4204, N4423, N4487, N4721, N4780, N5026, N5081, N5327, N5388, N5633, N5693, N5907, N5955, N1335, N1474, N1542, N1791, N1860, N2113, N2185, N2442, N2512, N2773, N2842, N3107, N3176, N3445, N3515, N3788, N3861, N4073, N4139, N4368, N4428, N4671, N4726, N4968, N5031, N5271, N5332, N5569, N5638, N5861, N5912, N1339, N1478, N1547, N1795, N1865, N2117, N2190, N2446, N2517, N2777, N2847, N3111, N3181, N3449, N3520, N3730, N3793, N4022, N4078, N4323, N4373, N4616, N4676, N4916, N4973, N5209, N5276, N5510, N5574, N5813, N5866, N1343, N1482, N1552, N1799, N1870, N2121, N2195, N2450, N2522, N2781, N2852, N3115, N3186, N3392, N3454, N3681, N3735, N3980, N4027, N4269, N4328, N4566, N4621, N4854, N4921, N5151, N5214, N5455, N5515, N5764, N5818, N1347, N1486, N1557, N1803, N1875, N2125, N2200, N2454, N2527, N2785, N2857, N3058, N3120, N3344, N3397, N3641, N3686, N3926, N3985, N4220, N4274, N4503, N4571, N4796, N4859, N5097, N5156, N5404, N5460, N5709, N5769, N1351, N1490, N1562, N1807, N1880, N2129, N2205, N2458, N2532, N2727, N2790, N3010, N3063, N3305, N3349, N3586, N3646, N3877, N3931, N4155, N4225, N4444, N4508, N4742, N4801, N5047, N5102, N5348, N5409, N5654, N5714, N1355, N1494, N1567, N1811, N1885, N2133, N2210, N2398, N2463, N2678, N2732, N2971, N3015, N3248, N3310, N3536, N3591, N3809, N3882, N4094, N4160, N4389, N4449, N4692, N4747, N4989, N5052, N5292, N5353, N5590, N5659, N1359, N1498, N1572, N1815, N1890, N2076, N2138, N2353, N2403, N2644, N2683, N2917, N2976, N3202, N3253, N3470, N3541, N3751, N3814, N4043, N4099, N4344, N4394, N4637, N4697, N4937, N4994, N5230, N5297, N5531, N5595, N1363, N1502, N1577, N1759, N1820, N2033, N2081, N2322, N2358, N2591, N2649, N2873, N2922, N3136, N3207, N3413, N3475, N3702, N3756, N4001, N4048, N4290, N4349, N4587, N4642, N4875, N4942, N5172, N5235, N5476, N5536, N1367, N1624, N1684, N1897, N1945, N2145, N2221, N2410, N2474, N2690, N2743, N2983, N3026, N3260, N3321, N3548, N3602, N3821, N3893, N4106, N4171, N4401, N4460, N4704, N4758, N5001, N5063, N5304, N5364, N5602, N5670, N1506, N1581, N1824, N1826, N1901, N2149, N2151, N2223, N2476, N2478, N2548, N2806, N2808, N2877, N3140, N3142, N3211, N3479, N3481, N3552, N3825, N3827, N3895, N4173, N4175, N4241, N4524, N4526, N4591, N4879, N4881, N4946, N5239, N5241, N5308, N5606, N5608, N5672, N5928, N5930, N5971, N6106, N6108, N6123, N1511, N1582, N1829, N1831, N1902, N2154, N2156, N2224, N2481, N2483, N2549, N2811, N2813, N2878, N3145, N3147, N3212, N3484, N3486, N3553, N3830, N3832, N3896, N4178, N4180, N4242, N4529, N4531, N4592, N4884, N4886, N4947, N5244, N5246, N5309, N5611, N5613, N5673, N5933, N5935, N5972, N6089, N6091, N6111, N1516, N1585, N1834, N1836, N1905, N2159, N2161, N2227, N2486, N2488, N2552, N2816, N2818, N2881, N3150, N3152, N3215, N3489, N3491, N3556, N3835, N3837, N3899, N4183, N4185, N4245, N4534, N4536, N4595, N4889, N4891, N4950, N5249, N5251, N5312, N5616, N5618, N5676, N5890, N5892, N5938, N6068, N6070, N6094, N1521, N1588, N1839, N1841, N1908, N2164, N2166, N2230, N2491, N2493, N2555, N2821, N2823, N2884, N3155, N3157, N3218, N3494, N3496, N3559, N3840, N3842, N3902, N4188, N4190, N4248, N4539, N4541, N4598, N4894, N4896, N4953, N5254, N5256, N5315, N5552, N5554, N5621, N5844, N5846, N5895, N6044, N6046, N6073, N1526, N1591, N1844, N1846, N1911, N2169, N2171, N2233, N2496, N2498, N2558, N2826, N2828, N2887, N3160, N3162, N3221, N3499, N3501, N3562, N3845, N3847, N3905, N4193, N4195, N4251, N4544, N4546, N4601, N4899, N4901, N4956, N5192, N5194, N5259, N5493, N5495, N5557, N5796, N5798, N5849, N6018, N6020, N6049, N1531, N1594, N1849, N1851, N1914, N2174, N2176, N2236, N2501, N2503, N2561, N2831, N2833, N2890, N3165, N3167, N3224, N3504, N3506, N3565, N3850, N3852, N3908, N4198, N4200, N4254, N4549, N4551, N4604, N4837, N4839, N4904, N5134, N5136, N5197, N5438, N5440, N5498, N5747, N5749, N5801, N5988, N5990, N6023, N1536, N1597, N1854, N1856, N1917, N2179, N2181, N2239, N2506, N2508, N2564, N2836, N2838, N2893, N3170, N3172, N3227, N3509, N3511, N3568, N3855, N3857, N3911, N4203, N4205, N4257, N4486, N4488, N4554, N4779, N4781, N4842, N5080, N5082, N5139, N5387, N5389, N5443, N5692, N5694, N5752, N5954, N5956, N5993, N1541, N1600, N1859, N1861, N1920, N2184, N2186, N2242, N2511, N2513, N2567, N2841, N2843, N2896, N3175, N3177, N3230, N3514, N3516, N3571, N3860, N3862, N3914, N4138, N4140, N4208, N4427, N4429, N4491, N4725, N4727, N4784, N5030, N5032, N5085, N5331, N5333, N5392, N5637, N5639, N5697, N5911, N5913, N5959, N1546, N1603, N1864, N1866, N1923, N2189, N2191, N2245, N2516, N2518, N2570, N2846, N2848, N2899, N3180, N3182, N3233, N3519, N3521, N3574, N3792, N3794, N3865, N4077, N4079, N4143, N4372, N4374, N4432, N4675, N4677, N4730, N4972, N4974, N5035, N5275, N5277, N5336, N5573, N5575, N5642, N5865, N5867, N5916, N1551, N1606, N1869, N1871, N1926, N2194, N2196, N2248, N2521, N2523, N2573, N2851, N2853, N2902, N3185, N3187, N3236, N3453, N3455, N3524, N3734, N3736, N3797, N4026, N4028, N4082, N4327, N4329, N4377, N4620, N4622, N4680, N4920, N4922, N4977, N5213, N5215, N5280, N5514, N5516, N5578, N5817, N5819, N5870, N1556, N1609, N1874, N1876, N1929, N2199, N2201, N2251, N2526, N2528, N2576, N2856, N2858, N2905, N3119, N3121, N3190, N3396, N3398, N3458, N3685, N3687, N3739, N3984, N3986, N4031, N4273, N4275, N4332, N4570, N4572, N4625, N4858, N4860, N4925, N5155, N5157, N5218, N5459, N5461, N5519, N5768, N5770, N5822, N1561, N1612, N1879, N1881, N1932, N2204, N2206, N2254, N2531, N2533, N2579, N2789, N2791, N2861, N3062, N3064, N3124, N3348, N3350, N3401, N3645, N3647, N3690, N3930, N3932, N3989, N4224, N4226, N4278, N4507, N4509, N4575, N4800, N4802, N4863, N5101, N5103, N5160, N5408, N5410, N5464, N5713, N5715, N5773, N1566, N1615, N1884, N1886, N1935, N2209, N2211, N2257, N2462, N2464, N2536, N2731, N2733, N2794, N3014, N3016, N3067, N3309, N3311, N3353, N3590, N3592, N3650, N3881, N3883, N3935, N4159, N4161, N4229, N4448, N4450, N4512, N4746, N4748, N4805, N5051, N5053, N5106, N5352, N5354, N5413, N5658, N5660, N5718, N1571, N1618, N1889, N1891, N1938, N2137, N2139, N2214, N2402, N2404, N2467, N2682, N2684, N2736, N2975, N2977, N3019, N3252, N3254, N3314, N3540, N3542, N3595, N3813, N3815, N3886, N4098, N4100, N4164, N4393, N4395, N4453, N4696, N4698, N4751, N4993, N4995, N5056, N5296, N5298, N5357, N5594, N5596, N5663, N1576, N1621, N1819, N1821, N1894, N2080, N2082, N2142, N2357, N2359, N2407, N2648, N2650, N2687, N2921, N2923, N2980, N3206, N3208, N3257, N3474, N3476, N3545, N3755, N3757, N3818, N4047, N4049, N4103, N4348, N4350, N4398, N4641, N4643, N4701, N4941, N4943, N4998, N5234, N5236, N5301, N5535, N5537, N5599, N1685, N1714, N1946, N2001, N2222, N2266, N2475, N2545, N2744, N2803, N3027, N3076, N3322, N3362, N3603, N3659, N3894, N3944, N4172, N4238, N4461, N4521, N4759, N4814, N5064, N5115, N5365, N5422, N5671, N6287, N5727, N1628, N1687, N1947, N2005, N2269, N2327, N2595, N2654, N2926, N2988, N3264, N3324, N3604, N3663, N3947, N4006, N4294, N4354, N4646, N4709, N5005, N5066, N5366, N5426, N5730, N5786, N6005, N6036, N6124, N6134, N1632, N1689, N1686, N1951, N2007, N2004, N2273, N2329, N2326, N2599, N2656, N2653, N2930, N2990, N2987, N3268, N3326, N3323, N3608, N3665, N3662, N3951, N4008, N4005, N4298, N4356, N4353, N4650, N4711, N4708, N5009, N5068, N5065, N5370, N5428, N5425, N5734, N5788, N5785, N5975, N6010, N6035, N6114, N6129, N6133, N1636, N1691, N1688, N1955, N2009, N2006, N2277, N2331, N2328, N2603, N2658, N2655, N2934, N2992, N2989, N3272, N3328, N3325, N3612, N3667, N3664, N3955, N4010, N4007, N4302, N4358, N4355, N4654, N4713, N4710, N5013, N5070, N5067, N5374, N5430, N5427, N5679, N5739, N5787, N5941, N5980, N6009, N6097, N6119, N6128, N1640, N1693, N1690, N1959, N2011, N2008, N2281, N2333, N2330, N2607, N2660, N2657, N2938, N2994, N2991, N3276, N3330, N3327, N3616, N3669, N3666, N3959, N4012, N4009, N4306, N4360, N4357, N4658, N4715, N4712, N5017, N5072, N5069, N5318, N5379, N5429, N5624, N5684, N5738, N5898, N5946, N5979, N6076, N6102, N6118, N1644, N1695, N1692, N1963, N2013, N2010, N2285, N2335, N2332, N2611, N2662, N2659, N2942, N2996, N2993, N3280, N3332, N3329, N3620, N3671, N3668, N3963, N4014, N4011, N4310, N4362, N4359, N4662, N4717, N4714, N4959, N5022, N5071, N5262, N5323, N5378, N5560, N5629, N5683, N5852, N5903, N5945, N6052, N6081, N6101, N1648, N1697, N1694, N1967, N2015, N2012, N2289, N2337, N2334, N2615, N2664, N2661, N2946, N2998, N2995, N3284, N3334, N3331, N3624, N3673, N3670, N3967, N4016, N4013, N4314, N4364, N4361, N4607, N4667, N4716, N4907, N4964, N5021, N5200, N5267, N5322, N5501, N5565, N5628, N5804, N5857, N5902, N6026, N6057, N6080, N1652, N1699, N1696, N1971, N2017, N2014, N2293, N2339, N2336, N2619, N2666, N2663, N2950, N3000, N2997, N3288, N3336, N3333, N3628, N3675, N3672, N3971, N4018, N4015, N4260, N4319, N4363, N4557, N4612, N4666, N4845, N4912, N4963, N5142, N5205, N5266, N5446, N5506, N5564, N5755, N5809, N5856, N5996, N6031, N6056, N1656, N1701, N1698, N1975, N2019, N2016, N2297, N2341, N2338, N2623, N2668, N2665, N2954, N3002, N2999, N3292, N3338, N3335, N3632, N3677, N3674, N3917, N3976, N4017, N4211, N4265, N4318, N4494, N4562, N4611, N4787, N4850, N4911, N5088, N5147, N5204, N5395, N5451, N5505, N5700, N5760, N5808, N5962, N6001, N6030, N1660, N1703, N1700, N1979, N2021, N2018, N2301, N2343, N2340, N2627, N2670, N2667, N2958, N3004, N3001, N3296, N3340, N3337, N3577, N3637, N3676, N3868, N3922, N3975, N4146, N4216, N4264, N4435, N4499, N4561, N4733, N4792, N4849, N5038, N5093, N5146, N5339, N5400, N5450, N5645, N5705, N5759, N5919, N5967, N6000, N1664, N1705, N1702, N1983, N2023, N2020, N2305, N2345, N2342, N2631, N2672, N2669, N2962, N3006, N3003, N3239, N3301, N3339, N3527, N3582, N3636, N3800, N3873, N3921, N4085, N4151, N4215, N4380, N4440, N4498, N4683, N4738, N4791, N4980, N5043, N5092, N5283, N5344, N5399, N5581, N5650, N5704, N5873, N5924, N5966, N1668, N1707, N1704, N1987, N2025, N2022, N2309, N2347, N2344, N2635, N2674, N2671, N2908, N2967, N3005, N3193, N3244, N3300, N3461, N3532, N3581, N3742, N3805, N3872, N4034, N4090, N4150, N4335, N4385, N4439, N4628, N4688, N4737, N4928, N4985, N5042, N5221, N5288, N5343, N5522, N5586, N5649, N5825, N5878, N5923, N1672, N1709, N1706, N1991, N2027, N2024, N2313, N2349, N2346, N2582, N2640, N2673, N2864, N2913, N2966, N3127, N3198, N3243, N3404, N3466, N3531, N3693, N3747, N3804, N3992, N4039, N4089, N4281, N4340, N4384, N4578, N4633, N4687, N4866, N4933, N4984, N5163, N5226, N5287, N5467, N5527, N5585, N5776, N5830, N5877, N1676, N1711, N1708, N1995, N2029, N2026, N2260, N2318, N2348, N2539, N2587, N2639, N2797, N2869, N2912, N3070, N3132, N3197, N3356, N3409, N3465, N3653, N3698, N3746, N3938, N3997, N4038, N4232, N4286, N4339, N4515, N4583, N4632, N4808, N4871, N4932, N5109, N5168, N5225, N5416, N5472, N5526, N5721, N5781, N5829, N1680, N1713, N1710, N1941, N2000, N2028, N2217, N2265, N2317, N2470, N2544, N2586, N2739, N2802, N2868, N3022, N3075, N3131, N3317, N3361, N3408, N3598, N3658, N3697, N3889, N3943, N3996, N4167, N4237, N4285, N4456, N4520, N4582, N4754, N4813, N4870, N5059, N5114, N5167, N5360, N5421, N5471, N5666, N5726, N5780, N1712, N1999, N2264, N2543, N2801, N3074, N3360, N3657, N3942, N4236, N4519, N4812, N5113, N5420, N5725, N6281, N6285, N1717, N2037, N2362, N2694, N3028, N3365, N3706, N4052, N4405, N4760, N5118, N5480, N5834, N6061, N6147, N6138, N1720, N2040, N2365, N2697, N3031, N3368, N3709, N4055, N4408, N4763, N5121, N5483, N5837, N6037, N6157, N6135, N1723, N2043, N2368, N2700, N3034, N3371, N3712, N4058, N4411, N4766, N5124, N5486, N5789, N6011, N6167, N6130, N1726, N2046, N2371, N2703, N3037, N3374, N3715, N4061, N4414, N4769, N5127, N5431, N5740, N5981, N6177, N6120, N1729, N2049, N2374, N2706, N3040, N3377, N3718, N4064, N4417, N4772, N5073, N5380, N5685, N5947, N6187, N6103, N1732, N2052, N2377, N2709, N3043, N3380, N3721, N4067, N4420, N4718, N5023, N5324, N5630, N5904, N6197, N6082, N1735, N2055, N2380, N2712, N3046, N3383, N3724, N4070, N4365, N4668, N4965, N5268, N5566, N5858, N6207, N6058, N1738, N2058, N2383, N2715, N3049, N3386, N3727, N4019, N4320, N4613, N4913, N5206, N5507, N5810, N6217, N6032, N1741, N2061, N2386, N2718, N3052, N3389, N3678, N3977, N4266, N4563, N4851, N5148, N5452, N5761, N6227, N6002, N1744, N2064, N2389, N2721, N3055, N3341, N3638, N3923, N4217, N4500, N4793, N5094, N5401, N5706, N6237, N5968, N1747, N2067, N2392, N2724, N3007, N3302, N3583, N3874, N4152, N4441, N4739, N5044, N5345, N5651, N6247, N5925, N1750, N2070, N2395, N2675, N2968, N3245, N3533, N3806, N4091, N4386, N4689, N4986, N5289, N5587, N6257, N5879, N1753, N2073, N2350, N2641, N2914, N3199, N3467, N3748, N4040, N4341, N4634, N4934, N5227, N5528, N6267, N5831, N1756, N2030, N2319, N2588, N2870, N3133, N3410, N3699, N3998, N4287, N4584, N4872, N5169, N5473, N6277, N5782, N6286, N6288, N6151, N6156, N6150, N6161, N6166, N6155, N6171, N6176, N6165, N6181, N6186, N6175, N6191, N6196, N6185, N6201, N6206, N6195, N6211, N6216, N6205, N6221, N6226, N6215, N6231, N6236, N6225, N6241, N6246, N6235, N6251, N6256, N6245, N6261, N6266, N6255, N6271, N6276, N6265, N6275, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280;
	assign N545 = ( N1 & N273 );
	assign N546 = ( N1 & N290 );
	assign N549 = ( N1 & N307 );
	assign N552 = ( N1 & N324 );
	assign N555 = ( N1 & N341 );
	assign N558 = ( N1 & N358 );
	assign N561 = ( N1 & N375 );
	assign N564 = ( N1 & N392 );
	assign N567 = ( N1 & N409 );
	assign N570 = ( N1 & N426 );
	assign N573 = ( N1 & N443 );
	assign N576 = ( N1 & N460 );
	assign N579 = ( N1 & N477 );
	assign N582 = ( N1 & N494 );
	assign N585 = ( N1 & N511 );
	assign N588 = ( N1 & N528 );
	assign N591 = ( N18 & N273 );
	assign N594 = ( N18 & N290 );
	assign N597 = ( N18 & N307 );
	assign N600 = ( N18 & N324 );
	assign N603 = ( N18 & N341 );
	assign N606 = ( N18 & N358 );
	assign N609 = ( N18 & N375 );
	assign N612 = ( N18 & N392 );
	assign N615 = ( N18 & N409 );
	assign N618 = ( N18 & N426 );
	assign N621 = ( N18 & N443 );
	assign N624 = ( N18 & N460 );
	assign N627 = ( N18 & N477 );
	assign N630 = ( N18 & N494 );
	assign N633 = ( N18 & N511 );
	assign N636 = ( N18 & N528 );
	assign N639 = ( N35 & N273 );
	assign N642 = ( N35 & N290 );
	assign N645 = ( N35 & N307 );
	assign N648 = ( N35 & N324 );
	assign N651 = ( N35 & N341 );
	assign N654 = ( N35 & N358 );
	assign N657 = ( N35 & N375 );
	assign N660 = ( N35 & N392 );
	assign N663 = ( N35 & N409 );
	assign N666 = ( N35 & N426 );
	assign N669 = ( N35 & N443 );
	assign N672 = ( N35 & N460 );
	assign N675 = ( N35 & N477 );
	assign N678 = ( N35 & N494 );
	assign N681 = ( N35 & N511 );
	assign N684 = ( N35 & N528 );
	assign N687 = ( N52 & N273 );
	assign N690 = ( N52 & N290 );
	assign N693 = ( N52 & N307 );
	assign N696 = ( N52 & N324 );
	assign N699 = ( N52 & N341 );
	assign N702 = ( N52 & N358 );
	assign N705 = ( N52 & N375 );
	assign N708 = ( N52 & N392 );
	assign N711 = ( N52 & N409 );
	assign N714 = ( N52 & N426 );
	assign N717 = ( N52 & N443 );
	assign N720 = ( N52 & N460 );
	assign N723 = ( N52 & N477 );
	assign N726 = ( N52 & N494 );
	assign N729 = ( N52 & N511 );
	assign N732 = ( N52 & N528 );
	assign N735 = ( N69 & N273 );
	assign N738 = ( N69 & N290 );
	assign N741 = ( N69 & N307 );
	assign N744 = ( N69 & N324 );
	assign N747 = ( N69 & N341 );
	assign N750 = ( N69 & N358 );
	assign N753 = ( N69 & N375 );
	assign N756 = ( N69 & N392 );
	assign N759 = ( N69 & N409 );
	assign N762 = ( N69 & N426 );
	assign N765 = ( N69 & N443 );
	assign N768 = ( N69 & N460 );
	assign N771 = ( N69 & N477 );
	assign N774 = ( N69 & N494 );
	assign N777 = ( N69 & N511 );
	assign N780 = ( N69 & N528 );
	assign N783 = ( N86 & N273 );
	assign N786 = ( N86 & N290 );
	assign N789 = ( N86 & N307 );
	assign N792 = ( N86 & N324 );
	assign N795 = ( N86 & N341 );
	assign N798 = ( N86 & N358 );
	assign N801 = ( N86 & N375 );
	assign N804 = ( N86 & N392 );
	assign N807 = ( N86 & N409 );
	assign N810 = ( N86 & N426 );
	assign N813 = ( N86 & N443 );
	assign N816 = ( N86 & N460 );
	assign N819 = ( N86 & N477 );
	assign N822 = ( N86 & N494 );
	assign N825 = ( N86 & N511 );
	assign N828 = ( N86 & N528 );
	assign N831 = ( N103 & N273 );
	assign N834 = ( N103 & N290 );
	assign N837 = ( N103 & N307 );
	assign N840 = ( N103 & N324 );
	assign N843 = ( N103 & N341 );
	assign N846 = ( N103 & N358 );
	assign N849 = ( N103 & N375 );
	assign N852 = ( N103 & N392 );
	assign N855 = ( N103 & N409 );
	assign N858 = ( N103 & N426 );
	assign N861 = ( N103 & N443 );
	assign N864 = ( N103 & N460 );
	assign N867 = ( N103 & N477 );
	assign N870 = ( N103 & N494 );
	assign N873 = ( N103 & N511 );
	assign N876 = ( N103 & N528 );
	assign N879 = ( N120 & N273 );
	assign N882 = ( N120 & N290 );
	assign N885 = ( N120 & N307 );
	assign N888 = ( N120 & N324 );
	assign N891 = ( N120 & N341 );
	assign N894 = ( N120 & N358 );
	assign N897 = ( N120 & N375 );
	assign N900 = ( N120 & N392 );
	assign N903 = ( N120 & N409 );
	assign N906 = ( N120 & N426 );
	assign N909 = ( N120 & N443 );
	assign N912 = ( N120 & N460 );
	assign N915 = ( N120 & N477 );
	assign N918 = ( N120 & N494 );
	assign N921 = ( N120 & N511 );
	assign N924 = ( N120 & N528 );
	assign N927 = ( N137 & N273 );
	assign N930 = ( N137 & N290 );
	assign N933 = ( N137 & N307 );
	assign N936 = ( N137 & N324 );
	assign N939 = ( N137 & N341 );
	assign N942 = ( N137 & N358 );
	assign N945 = ( N137 & N375 );
	assign N948 = ( N137 & N392 );
	assign N951 = ( N137 & N409 );
	assign N954 = ( N137 & N426 );
	assign N957 = ( N137 & N443 );
	assign N960 = ( N137 & N460 );
	assign N963 = ( N137 & N477 );
	assign N966 = ( N137 & N494 );
	assign N969 = ( N137 & N511 );
	assign N972 = ( N137 & N528 );
	assign N975 = ( N154 & N273 );
	assign N978 = ( N154 & N290 );
	assign N981 = ( N154 & N307 );
	assign N984 = ( N154 & N324 );
	assign N987 = ( N154 & N341 );
	assign N990 = ( N154 & N358 );
	assign N993 = ( N154 & N375 );
	assign N996 = ( N154 & N392 );
	assign N999 = ( N154 & N409 );
	assign N1002 = ( N154 & N426 );
	assign N1005 = ( N154 & N443 );
	assign N1008 = ( N154 & N460 );
	assign N1011 = ( N154 & N477 );
	assign N1014 = ( N154 & N494 );
	assign N1017 = ( N154 & N511 );
	assign N1020 = ( N154 & N528 );
	assign N1023 = ( N171 & N273 );
	assign N1026 = ( N171 & N290 );
	assign N1029 = ( N171 & N307 );
	assign N1032 = ( N171 & N324 );
	assign N1035 = ( N171 & N341 );
	assign N1038 = ( N171 & N358 );
	assign N1041 = ( N171 & N375 );
	assign N1044 = ( N171 & N392 );
	assign N1047 = ( N171 & N409 );
	assign N1050 = ( N171 & N426 );
	assign N1053 = ( N171 & N443 );
	assign N1056 = ( N171 & N460 );
	assign N1059 = ( N171 & N477 );
	assign N1062 = ( N171 & N494 );
	assign N1065 = ( N171 & N511 );
	assign N1068 = ( N171 & N528 );
	assign N1071 = ( N188 & N273 );
	assign N1074 = ( N188 & N290 );
	assign N1077 = ( N188 & N307 );
	assign N1080 = ( N188 & N324 );
	assign N1083 = ( N188 & N341 );
	assign N1086 = ( N188 & N358 );
	assign N1089 = ( N188 & N375 );
	assign N1092 = ( N188 & N392 );
	assign N1095 = ( N188 & N409 );
	assign N1098 = ( N188 & N426 );
	assign N1101 = ( N188 & N443 );
	assign N1104 = ( N188 & N460 );
	assign N1107 = ( N188 & N477 );
	assign N1110 = ( N188 & N494 );
	assign N1113 = ( N188 & N511 );
	assign N1116 = ( N188 & N528 );
	assign N1119 = ( N205 & N273 );
	assign N1122 = ( N205 & N290 );
	assign N1125 = ( N205 & N307 );
	assign N1128 = ( N205 & N324 );
	assign N1131 = ( N205 & N341 );
	assign N1134 = ( N205 & N358 );
	assign N1137 = ( N205 & N375 );
	assign N1140 = ( N205 & N392 );
	assign N1143 = ( N205 & N409 );
	assign N1146 = ( N205 & N426 );
	assign N1149 = ( N205 & N443 );
	assign N1152 = ( N205 & N460 );
	assign N1155 = ( N205 & N477 );
	assign N1158 = ( N205 & N494 );
	assign N1161 = ( N205 & N511 );
	assign N1164 = ( N205 & N528 );
	assign N1167 = ( N222 & N273 );
	assign N1170 = ( N222 & N290 );
	assign N1173 = ( N222 & N307 );
	assign N1176 = ( N222 & N324 );
	assign N1179 = ( N222 & N341 );
	assign N1182 = ( N222 & N358 );
	assign N1185 = ( N222 & N375 );
	assign N1188 = ( N222 & N392 );
	assign N1191 = ( N222 & N409 );
	assign N1194 = ( N222 & N426 );
	assign N1197 = ( N222 & N443 );
	assign N1200 = ( N222 & N460 );
	assign N1203 = ( N222 & N477 );
	assign N1206 = ( N222 & N494 );
	assign N1209 = ( N222 & N511 );
	assign N1212 = ( N222 & N528 );
	assign N1215 = ( N239 & N273 );
	assign N1218 = ( N239 & N290 );
	assign N1221 = ( N239 & N307 );
	assign N1224 = ( N239 & N324 );
	assign N1227 = ( N239 & N341 );
	assign N1230 = ( N239 & N358 );
	assign N1233 = ( N239 & N375 );
	assign N1236 = ( N239 & N392 );
	assign N1239 = ( N239 & N409 );
	assign N1242 = ( N239 & N426 );
	assign N1245 = ( N239 & N443 );
	assign N1248 = ( N239 & N460 );
	assign N1251 = ( N239 & N477 );
	assign N1254 = ( N239 & N494 );
	assign N1257 = ( N239 & N511 );
	assign N1260 = ( N239 & N528 );
	assign N1263 = ( N256 & N273 );
	assign N1266 = ( N256 & N290 );
	assign N1269 = ( N256 & N307 );
	assign N1272 = ( N256 & N324 );
	assign N1275 = ( N256 & N341 );
	assign N1278 = ( N256 & N358 );
	assign N1281 = ( N256 & N375 );
	assign N1284 = ( N256 & N392 );
	assign N1287 = ( N256 & N409 );
	assign N1290 = ( N256 & N426 );
	assign N1293 = ( N256 & N443 );
	assign N1296 = ( N256 & N460 );
	assign N1299 = ( N256 & N477 );
	assign N1302 = ( N256 & N494 );
	assign N1305 = ( N256 & N511 );
	assign N1308 = ( N256 & N528 );
	assign N1446 = ~( N1311 | N546 );
	assign N1507 = ~( N1446 | N546 );
	assign N1763 = ~( N1717 | N549 );
	assign N1825 = ~( N1763 | N549 );
	assign N2085 = ~( N2037 | N552 );
	assign N2150 = ~( N2085 | N552 );
	assign N2414 = ~( N2362 | N555 );
	assign N2477 = ~( N2414 | N555 );
	assign N2745 = ~( N2694 | N558 );
	assign N2807 = ~( N2745 | N558 );
	assign N3079 = ~( N3028 | N561 );
	assign N3141 = ~( N3079 | N561 );
	assign N3417 = ~( N3365 | N564 );
	assign N3480 = ~( N3417 | N564 );
	assign N3760 = ~( N3706 | N567 );
	assign N3826 = ~( N3760 | N567 );
	assign N4110 = ~( N4052 | N570 );
	assign N4174 = ~( N4110 | N570 );
	assign N4462 = ~( N4405 | N573 );
	assign N4525 = ~( N4462 | N573 );
	assign N4817 = ~( N4760 | N576 );
	assign N4880 = ~( N4817 | N576 );
	assign N5176 = ~( N5118 | N579 );
	assign N5240 = ~( N5176 | N579 );
	assign N5540 = ~( N5480 | N582 );
	assign N5607 = ~( N5540 | N582 );
	assign N5882 = ~( N5834 | N585 );
	assign N5929 = ~( N5882 | N585 );
	assign N6085 = ~( N6061 | N588 );
	assign N6107 = ~( N6085 | N588 );
	assign N1311 = ~N591;
	assign N1450 = ~( N1315 | N594 );
	assign N1512 = ~( N1450 | N594 );
	assign N1767 = ~( N1720 | N597 );
	assign N1830 = ~( N1767 | N597 );
	assign N2089 = ~( N2040 | N600 );
	assign N2155 = ~( N2089 | N600 );
	assign N2418 = ~( N2365 | N603 );
	assign N2482 = ~( N2418 | N603 );
	assign N2749 = ~( N2697 | N606 );
	assign N2812 = ~( N2749 | N606 );
	assign N3083 = ~( N3031 | N609 );
	assign N3146 = ~( N3083 | N609 );
	assign N3421 = ~( N3368 | N612 );
	assign N3485 = ~( N3421 | N612 );
	assign N3764 = ~( N3709 | N615 );
	assign N3831 = ~( N3764 | N615 );
	assign N4114 = ~( N4055 | N618 );
	assign N4179 = ~( N4114 | N618 );
	assign N4466 = ~( N4408 | N621 );
	assign N4530 = ~( N4466 | N621 );
	assign N4821 = ~( N4763 | N624 );
	assign N4885 = ~( N4821 | N624 );
	assign N5180 = ~( N5121 | N627 );
	assign N5245 = ~( N5180 | N627 );
	assign N5544 = ~( N5483 | N630 );
	assign N5612 = ~( N5544 | N630 );
	assign N5886 = ~( N5837 | N633 );
	assign N5934 = ~( N5886 | N633 );
	assign N6064 = ~( N6037 | N636 );
	assign N6090 = ~( N6064 | N636 );
	assign N1315 = ~N639;
	assign N1454 = ~( N1319 | N642 );
	assign N1517 = ~( N1454 | N642 );
	assign N1771 = ~( N1723 | N645 );
	assign N1835 = ~( N1771 | N645 );
	assign N2093 = ~( N2043 | N648 );
	assign N2160 = ~( N2093 | N648 );
	assign N2422 = ~( N2368 | N651 );
	assign N2487 = ~( N2422 | N651 );
	assign N2753 = ~( N2700 | N654 );
	assign N2817 = ~( N2753 | N654 );
	assign N3087 = ~( N3034 | N657 );
	assign N3151 = ~( N3087 | N657 );
	assign N3425 = ~( N3371 | N660 );
	assign N3490 = ~( N3425 | N660 );
	assign N3768 = ~( N3712 | N663 );
	assign N3836 = ~( N3768 | N663 );
	assign N4118 = ~( N4058 | N666 );
	assign N4184 = ~( N4118 | N666 );
	assign N4470 = ~( N4411 | N669 );
	assign N4535 = ~( N4470 | N669 );
	assign N4825 = ~( N4766 | N672 );
	assign N4890 = ~( N4825 | N672 );
	assign N5184 = ~( N5124 | N675 );
	assign N5250 = ~( N5184 | N675 );
	assign N5548 = ~( N5486 | N678 );
	assign N5617 = ~( N5548 | N678 );
	assign N5840 = ~( N5789 | N681 );
	assign N5891 = ~( N5840 | N681 );
	assign N6040 = ~( N6011 | N684 );
	assign N6069 = ~( N6040 | N684 );
	assign N1319 = ~N687;
	assign N1458 = ~( N1323 | N690 );
	assign N1522 = ~( N1458 | N690 );
	assign N1775 = ~( N1726 | N693 );
	assign N1840 = ~( N1775 | N693 );
	assign N2097 = ~( N2046 | N696 );
	assign N2165 = ~( N2097 | N696 );
	assign N2426 = ~( N2371 | N699 );
	assign N2492 = ~( N2426 | N699 );
	assign N2757 = ~( N2703 | N702 );
	assign N2822 = ~( N2757 | N702 );
	assign N3091 = ~( N3037 | N705 );
	assign N3156 = ~( N3091 | N705 );
	assign N3429 = ~( N3374 | N708 );
	assign N3495 = ~( N3429 | N708 );
	assign N3772 = ~( N3715 | N711 );
	assign N3841 = ~( N3772 | N711 );
	assign N4122 = ~( N4061 | N714 );
	assign N4189 = ~( N4122 | N714 );
	assign N4474 = ~( N4414 | N717 );
	assign N4540 = ~( N4474 | N717 );
	assign N4829 = ~( N4769 | N720 );
	assign N4895 = ~( N4829 | N720 );
	assign N5188 = ~( N5127 | N723 );
	assign N5255 = ~( N5188 | N723 );
	assign N5489 = ~( N5431 | N726 );
	assign N5553 = ~( N5489 | N726 );
	assign N5792 = ~( N5740 | N729 );
	assign N5845 = ~( N5792 | N729 );
	assign N6014 = ~( N5981 | N732 );
	assign N6045 = ~( N6014 | N732 );
	assign N1323 = ~N735;
	assign N1462 = ~( N1327 | N738 );
	assign N1527 = ~( N1462 | N738 );
	assign N1779 = ~( N1729 | N741 );
	assign N1845 = ~( N1779 | N741 );
	assign N2101 = ~( N2049 | N744 );
	assign N2170 = ~( N2101 | N744 );
	assign N2430 = ~( N2374 | N747 );
	assign N2497 = ~( N2430 | N747 );
	assign N2761 = ~( N2706 | N750 );
	assign N2827 = ~( N2761 | N750 );
	assign N3095 = ~( N3040 | N753 );
	assign N3161 = ~( N3095 | N753 );
	assign N3433 = ~( N3377 | N756 );
	assign N3500 = ~( N3433 | N756 );
	assign N3776 = ~( N3718 | N759 );
	assign N3846 = ~( N3776 | N759 );
	assign N4126 = ~( N4064 | N762 );
	assign N4194 = ~( N4126 | N762 );
	assign N4478 = ~( N4417 | N765 );
	assign N4545 = ~( N4478 | N765 );
	assign N4833 = ~( N4772 | N768 );
	assign N4900 = ~( N4833 | N768 );
	assign N5130 = ~( N5073 | N771 );
	assign N5193 = ~( N5130 | N771 );
	assign N5434 = ~( N5380 | N774 );
	assign N5494 = ~( N5434 | N774 );
	assign N5743 = ~( N5685 | N777 );
	assign N5797 = ~( N5743 | N777 );
	assign N5984 = ~( N5947 | N780 );
	assign N6019 = ~( N5984 | N780 );
	assign N1327 = ~N783;
	assign N1466 = ~( N1331 | N786 );
	assign N1532 = ~( N1466 | N786 );
	assign N1783 = ~( N1732 | N789 );
	assign N1850 = ~( N1783 | N789 );
	assign N2105 = ~( N2052 | N792 );
	assign N2175 = ~( N2105 | N792 );
	assign N2434 = ~( N2377 | N795 );
	assign N2502 = ~( N2434 | N795 );
	assign N2765 = ~( N2709 | N798 );
	assign N2832 = ~( N2765 | N798 );
	assign N3099 = ~( N3043 | N801 );
	assign N3166 = ~( N3099 | N801 );
	assign N3437 = ~( N3380 | N804 );
	assign N3505 = ~( N3437 | N804 );
	assign N3780 = ~( N3721 | N807 );
	assign N3851 = ~( N3780 | N807 );
	assign N4130 = ~( N4067 | N810 );
	assign N4199 = ~( N4130 | N810 );
	assign N4482 = ~( N4420 | N813 );
	assign N4550 = ~( N4482 | N813 );
	assign N4775 = ~( N4718 | N816 );
	assign N4838 = ~( N4775 | N816 );
	assign N5076 = ~( N5023 | N819 );
	assign N5135 = ~( N5076 | N819 );
	assign N5383 = ~( N5324 | N822 );
	assign N5439 = ~( N5383 | N822 );
	assign N5688 = ~( N5630 | N825 );
	assign N5748 = ~( N5688 | N825 );
	assign N5950 = ~( N5904 | N828 );
	assign N5989 = ~( N5950 | N828 );
	assign N1331 = ~N831;
	assign N1470 = ~( N1335 | N834 );
	assign N1537 = ~( N1470 | N834 );
	assign N1787 = ~( N1735 | N837 );
	assign N1855 = ~( N1787 | N837 );
	assign N2109 = ~( N2055 | N840 );
	assign N2180 = ~( N2109 | N840 );
	assign N2438 = ~( N2380 | N843 );
	assign N2507 = ~( N2438 | N843 );
	assign N2769 = ~( N2712 | N846 );
	assign N2837 = ~( N2769 | N846 );
	assign N3103 = ~( N3046 | N849 );
	assign N3171 = ~( N3103 | N849 );
	assign N3441 = ~( N3383 | N852 );
	assign N3510 = ~( N3441 | N852 );
	assign N3784 = ~( N3724 | N855 );
	assign N3856 = ~( N3784 | N855 );
	assign N4134 = ~( N4070 | N858 );
	assign N4204 = ~( N4134 | N858 );
	assign N4423 = ~( N4365 | N861 );
	assign N4487 = ~( N4423 | N861 );
	assign N4721 = ~( N4668 | N864 );
	assign N4780 = ~( N4721 | N864 );
	assign N5026 = ~( N4965 | N867 );
	assign N5081 = ~( N5026 | N867 );
	assign N5327 = ~( N5268 | N870 );
	assign N5388 = ~( N5327 | N870 );
	assign N5633 = ~( N5566 | N873 );
	assign N5693 = ~( N5633 | N873 );
	assign N5907 = ~( N5858 | N876 );
	assign N5955 = ~( N5907 | N876 );
	assign N1335 = ~N879;
	assign N1474 = ~( N1339 | N882 );
	assign N1542 = ~( N1474 | N882 );
	assign N1791 = ~( N1738 | N885 );
	assign N1860 = ~( N1791 | N885 );
	assign N2113 = ~( N2058 | N888 );
	assign N2185 = ~( N2113 | N888 );
	assign N2442 = ~( N2383 | N891 );
	assign N2512 = ~( N2442 | N891 );
	assign N2773 = ~( N2715 | N894 );
	assign N2842 = ~( N2773 | N894 );
	assign N3107 = ~( N3049 | N897 );
	assign N3176 = ~( N3107 | N897 );
	assign N3445 = ~( N3386 | N900 );
	assign N3515 = ~( N3445 | N900 );
	assign N3788 = ~( N3727 | N903 );
	assign N3861 = ~( N3788 | N903 );
	assign N4073 = ~( N4019 | N906 );
	assign N4139 = ~( N4073 | N906 );
	assign N4368 = ~( N4320 | N909 );
	assign N4428 = ~( N4368 | N909 );
	assign N4671 = ~( N4613 | N912 );
	assign N4726 = ~( N4671 | N912 );
	assign N4968 = ~( N4913 | N915 );
	assign N5031 = ~( N4968 | N915 );
	assign N5271 = ~( N5206 | N918 );
	assign N5332 = ~( N5271 | N918 );
	assign N5569 = ~( N5507 | N921 );
	assign N5638 = ~( N5569 | N921 );
	assign N5861 = ~( N5810 | N924 );
	assign N5912 = ~( N5861 | N924 );
	assign N1339 = ~N927;
	assign N1478 = ~( N1343 | N930 );
	assign N1547 = ~( N1478 | N930 );
	assign N1795 = ~( N1741 | N933 );
	assign N1865 = ~( N1795 | N933 );
	assign N2117 = ~( N2061 | N936 );
	assign N2190 = ~( N2117 | N936 );
	assign N2446 = ~( N2386 | N939 );
	assign N2517 = ~( N2446 | N939 );
	assign N2777 = ~( N2718 | N942 );
	assign N2847 = ~( N2777 | N942 );
	assign N3111 = ~( N3052 | N945 );
	assign N3181 = ~( N3111 | N945 );
	assign N3449 = ~( N3389 | N948 );
	assign N3520 = ~( N3449 | N948 );
	assign N3730 = ~( N3678 | N951 );
	assign N3793 = ~( N3730 | N951 );
	assign N4022 = ~( N3977 | N954 );
	assign N4078 = ~( N4022 | N954 );
	assign N4323 = ~( N4266 | N957 );
	assign N4373 = ~( N4323 | N957 );
	assign N4616 = ~( N4563 | N960 );
	assign N4676 = ~( N4616 | N960 );
	assign N4916 = ~( N4851 | N963 );
	assign N4973 = ~( N4916 | N963 );
	assign N5209 = ~( N5148 | N966 );
	assign N5276 = ~( N5209 | N966 );
	assign N5510 = ~( N5452 | N969 );
	assign N5574 = ~( N5510 | N969 );
	assign N5813 = ~( N5761 | N972 );
	assign N5866 = ~( N5813 | N972 );
	assign N1343 = ~N975;
	assign N1482 = ~( N1347 | N978 );
	assign N1552 = ~( N1482 | N978 );
	assign N1799 = ~( N1744 | N981 );
	assign N1870 = ~( N1799 | N981 );
	assign N2121 = ~( N2064 | N984 );
	assign N2195 = ~( N2121 | N984 );
	assign N2450 = ~( N2389 | N987 );
	assign N2522 = ~( N2450 | N987 );
	assign N2781 = ~( N2721 | N990 );
	assign N2852 = ~( N2781 | N990 );
	assign N3115 = ~( N3055 | N993 );
	assign N3186 = ~( N3115 | N993 );
	assign N3392 = ~( N3341 | N996 );
	assign N3454 = ~( N3392 | N996 );
	assign N3681 = ~( N3638 | N999 );
	assign N3735 = ~( N3681 | N999 );
	assign N3980 = ~( N3923 | N1002 );
	assign N4027 = ~( N3980 | N1002 );
	assign N4269 = ~( N4217 | N1005 );
	assign N4328 = ~( N4269 | N1005 );
	assign N4566 = ~( N4500 | N1008 );
	assign N4621 = ~( N4566 | N1008 );
	assign N4854 = ~( N4793 | N1011 );
	assign N4921 = ~( N4854 | N1011 );
	assign N5151 = ~( N5094 | N1014 );
	assign N5214 = ~( N5151 | N1014 );
	assign N5455 = ~( N5401 | N1017 );
	assign N5515 = ~( N5455 | N1017 );
	assign N5764 = ~( N5706 | N1020 );
	assign N5818 = ~( N5764 | N1020 );
	assign N1347 = ~N1023;
	assign N1486 = ~( N1351 | N1026 );
	assign N1557 = ~( N1486 | N1026 );
	assign N1803 = ~( N1747 | N1029 );
	assign N1875 = ~( N1803 | N1029 );
	assign N2125 = ~( N2067 | N1032 );
	assign N2200 = ~( N2125 | N1032 );
	assign N2454 = ~( N2392 | N1035 );
	assign N2527 = ~( N2454 | N1035 );
	assign N2785 = ~( N2724 | N1038 );
	assign N2857 = ~( N2785 | N1038 );
	assign N3058 = ~( N3007 | N1041 );
	assign N3120 = ~( N3058 | N1041 );
	assign N3344 = ~( N3302 | N1044 );
	assign N3397 = ~( N3344 | N1044 );
	assign N3641 = ~( N3583 | N1047 );
	assign N3686 = ~( N3641 | N1047 );
	assign N3926 = ~( N3874 | N1050 );
	assign N3985 = ~( N3926 | N1050 );
	assign N4220 = ~( N4152 | N1053 );
	assign N4274 = ~( N4220 | N1053 );
	assign N4503 = ~( N4441 | N1056 );
	assign N4571 = ~( N4503 | N1056 );
	assign N4796 = ~( N4739 | N1059 );
	assign N4859 = ~( N4796 | N1059 );
	assign N5097 = ~( N5044 | N1062 );
	assign N5156 = ~( N5097 | N1062 );
	assign N5404 = ~( N5345 | N1065 );
	assign N5460 = ~( N5404 | N1065 );
	assign N5709 = ~( N5651 | N1068 );
	assign N5769 = ~( N5709 | N1068 );
	assign N1351 = ~N1071;
	assign N1490 = ~( N1355 | N1074 );
	assign N1562 = ~( N1490 | N1074 );
	assign N1807 = ~( N1750 | N1077 );
	assign N1880 = ~( N1807 | N1077 );
	assign N2129 = ~( N2070 | N1080 );
	assign N2205 = ~( N2129 | N1080 );
	assign N2458 = ~( N2395 | N1083 );
	assign N2532 = ~( N2458 | N1083 );
	assign N2727 = ~( N2675 | N1086 );
	assign N2790 = ~( N2727 | N1086 );
	assign N3010 = ~( N2968 | N1089 );
	assign N3063 = ~( N3010 | N1089 );
	assign N3305 = ~( N3245 | N1092 );
	assign N3349 = ~( N3305 | N1092 );
	assign N3586 = ~( N3533 | N1095 );
	assign N3646 = ~( N3586 | N1095 );
	assign N3877 = ~( N3806 | N1098 );
	assign N3931 = ~( N3877 | N1098 );
	assign N4155 = ~( N4091 | N1101 );
	assign N4225 = ~( N4155 | N1101 );
	assign N4444 = ~( N4386 | N1104 );
	assign N4508 = ~( N4444 | N1104 );
	assign N4742 = ~( N4689 | N1107 );
	assign N4801 = ~( N4742 | N1107 );
	assign N5047 = ~( N4986 | N1110 );
	assign N5102 = ~( N5047 | N1110 );
	assign N5348 = ~( N5289 | N1113 );
	assign N5409 = ~( N5348 | N1113 );
	assign N5654 = ~( N5587 | N1116 );
	assign N5714 = ~( N5654 | N1116 );
	assign N1355 = ~N1119;
	assign N1494 = ~( N1359 | N1122 );
	assign N1567 = ~( N1494 | N1122 );
	assign N1811 = ~( N1753 | N1125 );
	assign N1885 = ~( N1811 | N1125 );
	assign N2133 = ~( N2073 | N1128 );
	assign N2210 = ~( N2133 | N1128 );
	assign N2398 = ~( N2350 | N1131 );
	assign N2463 = ~( N2398 | N1131 );
	assign N2678 = ~( N2641 | N1134 );
	assign N2732 = ~( N2678 | N1134 );
	assign N2971 = ~( N2914 | N1137 );
	assign N3015 = ~( N2971 | N1137 );
	assign N3248 = ~( N3199 | N1140 );
	assign N3310 = ~( N3248 | N1140 );
	assign N3536 = ~( N3467 | N1143 );
	assign N3591 = ~( N3536 | N1143 );
	assign N3809 = ~( N3748 | N1146 );
	assign N3882 = ~( N3809 | N1146 );
	assign N4094 = ~( N4040 | N1149 );
	assign N4160 = ~( N4094 | N1149 );
	assign N4389 = ~( N4341 | N1152 );
	assign N4449 = ~( N4389 | N1152 );
	assign N4692 = ~( N4634 | N1155 );
	assign N4747 = ~( N4692 | N1155 );
	assign N4989 = ~( N4934 | N1158 );
	assign N5052 = ~( N4989 | N1158 );
	assign N5292 = ~( N5227 | N1161 );
	assign N5353 = ~( N5292 | N1161 );
	assign N5590 = ~( N5528 | N1164 );
	assign N5659 = ~( N5590 | N1164 );
	assign N1359 = ~N1167;
	assign N1498 = ~( N1363 | N1170 );
	assign N1572 = ~( N1498 | N1170 );
	assign N1815 = ~( N1756 | N1173 );
	assign N1890 = ~( N1815 | N1173 );
	assign N2076 = ~( N2030 | N1176 );
	assign N2138 = ~( N2076 | N1176 );
	assign N2353 = ~( N2319 | N1179 );
	assign N2403 = ~( N2353 | N1179 );
	assign N2644 = ~( N2588 | N1182 );
	assign N2683 = ~( N2644 | N1182 );
	assign N2917 = ~( N2870 | N1185 );
	assign N2976 = ~( N2917 | N1185 );
	assign N3202 = ~( N3133 | N1188 );
	assign N3253 = ~( N3202 | N1188 );
	assign N3470 = ~( N3410 | N1191 );
	assign N3541 = ~( N3470 | N1191 );
	assign N3751 = ~( N3699 | N1194 );
	assign N3814 = ~( N3751 | N1194 );
	assign N4043 = ~( N3998 | N1197 );
	assign N4099 = ~( N4043 | N1197 );
	assign N4344 = ~( N4287 | N1200 );
	assign N4394 = ~( N4344 | N1200 );
	assign N4637 = ~( N4584 | N1203 );
	assign N4697 = ~( N4637 | N1203 );
	assign N4937 = ~( N4872 | N1206 );
	assign N4994 = ~( N4937 | N1206 );
	assign N5230 = ~( N5169 | N1209 );
	assign N5297 = ~( N5230 | N1209 );
	assign N5531 = ~( N5473 | N1212 );
	assign N5595 = ~( N5531 | N1212 );
	assign N1363 = ~N1215;
	assign N1502 = ~( N1367 | N1218 );
	assign N1577 = ~( N1502 | N1218 );
	assign N1759 = ~( N1714 | N1221 );
	assign N1820 = ~( N1759 | N1221 );
	assign N2033 = ~( N2001 | N1224 );
	assign N2081 = ~( N2033 | N1224 );
	assign N2322 = ~( N2266 | N1227 );
	assign N2358 = ~( N2322 | N1227 );
	assign N2591 = ~( N2545 | N1230 );
	assign N2649 = ~( N2591 | N1230 );
	assign N2873 = ~( N2803 | N1233 );
	assign N2922 = ~( N2873 | N1233 );
	assign N3136 = ~( N3076 | N1236 );
	assign N3207 = ~( N3136 | N1236 );
	assign N3413 = ~( N3362 | N1239 );
	assign N3475 = ~( N3413 | N1239 );
	assign N3702 = ~( N3659 | N1242 );
	assign N3756 = ~( N3702 | N1242 );
	assign N4001 = ~( N3944 | N1245 );
	assign N4048 = ~( N4001 | N1245 );
	assign N4290 = ~( N4238 | N1248 );
	assign N4349 = ~( N4290 | N1248 );
	assign N4587 = ~( N4521 | N1251 );
	assign N4642 = ~( N4587 | N1251 );
	assign N4875 = ~( N4814 | N1254 );
	assign N4942 = ~( N4875 | N1254 );
	assign N5172 = ~( N5115 | N1257 );
	assign N5235 = ~( N5172 | N1257 );
	assign N5476 = ~( N5422 | N1260 );
	assign N5536 = ~( N5476 | N1260 );
	assign N1367 = ~N1263;
	assign N1624 = ~( N1266 | N1576 );
	assign N1684 = ~( N1266 | N1624 );
	assign N1897 = ~( N1269 | N1821 );
	assign N1945 = ~( N1269 | N1897 );
	assign N2145 = ~( N1272 | N2082 );
	assign N2221 = ~( N1272 | N2145 );
	assign N2410 = ~( N1275 | N2359 );
	assign N2474 = ~( N1275 | N2410 );
	assign N2690 = ~( N1278 | N2650 );
	assign N2743 = ~( N1278 | N2690 );
	assign N2983 = ~( N1281 | N2923 );
	assign N3026 = ~( N1281 | N2983 );
	assign N3260 = ~( N1284 | N3208 );
	assign N3321 = ~( N1284 | N3260 );
	assign N3548 = ~( N1287 | N3476 );
	assign N3602 = ~( N1287 | N3548 );
	assign N3821 = ~( N1290 | N3757 );
	assign N3893 = ~( N1290 | N3821 );
	assign N4106 = ~( N1293 | N4049 );
	assign N4171 = ~( N1293 | N4106 );
	assign N4401 = ~( N1296 | N4350 );
	assign N4460 = ~( N1296 | N4401 );
	assign N4704 = ~( N1299 | N4643 );
	assign N4758 = ~( N1299 | N4704 );
	assign N5001 = ~( N1302 | N4943 );
	assign N5063 = ~( N1302 | N5001 );
	assign N5304 = ~( N1305 | N5236 );
	assign N5364 = ~( N1305 | N5304 );
	assign N5602 = ~( N1308 | N5537 );
	assign N5670 = ~( N1308 | N5602 );
	assign N1506 = ~( N1311 | N1446 );
	assign N1581 = ~( N1506 | N1507 );
	assign N1824 = ~( N1717 | N1763 );
	assign N1826 = ~( N1628 | N1763 );
	assign N1901 = ~( N1824 | N1825 );
	assign N2149 = ~( N2037 | N2085 );
	assign N2151 = ~( N1947 | N2085 );
	assign N2223 = ~( N2149 | N2150 );
	assign N2476 = ~( N2362 | N2414 );
	assign N2478 = ~( N2269 | N2414 );
	assign N2548 = ~( N2476 | N2477 );
	assign N2806 = ~( N2694 | N2745 );
	assign N2808 = ~( N2595 | N2745 );
	assign N2877 = ~( N2806 | N2807 );
	assign N3140 = ~( N3028 | N3079 );
	assign N3142 = ~( N2926 | N3079 );
	assign N3211 = ~( N3140 | N3141 );
	assign N3479 = ~( N3365 | N3417 );
	assign N3481 = ~( N3264 | N3417 );
	assign N3552 = ~( N3479 | N3480 );
	assign N3825 = ~( N3706 | N3760 );
	assign N3827 = ~( N3604 | N3760 );
	assign N3895 = ~( N3825 | N3826 );
	assign N4173 = ~( N4052 | N4110 );
	assign N4175 = ~( N3947 | N4110 );
	assign N4241 = ~( N4173 | N4174 );
	assign N4524 = ~( N4405 | N4462 );
	assign N4526 = ~( N4294 | N4462 );
	assign N4591 = ~( N4524 | N4525 );
	assign N4879 = ~( N4760 | N4817 );
	assign N4881 = ~( N4646 | N4817 );
	assign N4946 = ~( N4879 | N4880 );
	assign N5239 = ~( N5118 | N5176 );
	assign N5241 = ~( N5005 | N5176 );
	assign N5308 = ~( N5239 | N5240 );
	assign N5606 = ~( N5480 | N5540 );
	assign N5608 = ~( N5366 | N5540 );
	assign N5672 = ~( N5606 | N5607 );
	assign N5928 = ~( N5834 | N5882 );
	assign N5930 = ~( N5730 | N5882 );
	assign N5971 = ~( N5928 | N5929 );
	assign N6106 = ~( N6061 | N6085 );
	assign N6108 = ~( N6005 | N6085 );
	assign N6123 = ~( N6106 | N6107 );
	assign N1511 = ~( N1315 | N1450 );
	assign N1582 = ~( N1511 | N1512 );
	assign N1829 = ~( N1720 | N1767 );
	assign N1831 = ~( N1632 | N1767 );
	assign N1902 = ~( N1829 | N1830 );
	assign N2154 = ~( N2040 | N2089 );
	assign N2156 = ~( N1951 | N2089 );
	assign N2224 = ~( N2154 | N2155 );
	assign N2481 = ~( N2365 | N2418 );
	assign N2483 = ~( N2273 | N2418 );
	assign N2549 = ~( N2481 | N2482 );
	assign N2811 = ~( N2697 | N2749 );
	assign N2813 = ~( N2599 | N2749 );
	assign N2878 = ~( N2811 | N2812 );
	assign N3145 = ~( N3031 | N3083 );
	assign N3147 = ~( N2930 | N3083 );
	assign N3212 = ~( N3145 | N3146 );
	assign N3484 = ~( N3368 | N3421 );
	assign N3486 = ~( N3268 | N3421 );
	assign N3553 = ~( N3484 | N3485 );
	assign N3830 = ~( N3709 | N3764 );
	assign N3832 = ~( N3608 | N3764 );
	assign N3896 = ~( N3830 | N3831 );
	assign N4178 = ~( N4055 | N4114 );
	assign N4180 = ~( N3951 | N4114 );
	assign N4242 = ~( N4178 | N4179 );
	assign N4529 = ~( N4408 | N4466 );
	assign N4531 = ~( N4298 | N4466 );
	assign N4592 = ~( N4529 | N4530 );
	assign N4884 = ~( N4763 | N4821 );
	assign N4886 = ~( N4650 | N4821 );
	assign N4947 = ~( N4884 | N4885 );
	assign N5244 = ~( N5121 | N5180 );
	assign N5246 = ~( N5009 | N5180 );
	assign N5309 = ~( N5244 | N5245 );
	assign N5611 = ~( N5483 | N5544 );
	assign N5613 = ~( N5370 | N5544 );
	assign N5673 = ~( N5611 | N5612 );
	assign N5933 = ~( N5837 | N5886 );
	assign N5935 = ~( N5734 | N5886 );
	assign N5972 = ~( N5933 | N5934 );
	assign N6089 = ~( N6037 | N6064 );
	assign N6091 = ~( N5975 | N6064 );
	assign N6111 = ~( N6089 | N6090 );
	assign N1516 = ~( N1319 | N1454 );
	assign N1585 = ~( N1516 | N1517 );
	assign N1834 = ~( N1723 | N1771 );
	assign N1836 = ~( N1636 | N1771 );
	assign N1905 = ~( N1834 | N1835 );
	assign N2159 = ~( N2043 | N2093 );
	assign N2161 = ~( N1955 | N2093 );
	assign N2227 = ~( N2159 | N2160 );
	assign N2486 = ~( N2368 | N2422 );
	assign N2488 = ~( N2277 | N2422 );
	assign N2552 = ~( N2486 | N2487 );
	assign N2816 = ~( N2700 | N2753 );
	assign N2818 = ~( N2603 | N2753 );
	assign N2881 = ~( N2816 | N2817 );
	assign N3150 = ~( N3034 | N3087 );
	assign N3152 = ~( N2934 | N3087 );
	assign N3215 = ~( N3150 | N3151 );
	assign N3489 = ~( N3371 | N3425 );
	assign N3491 = ~( N3272 | N3425 );
	assign N3556 = ~( N3489 | N3490 );
	assign N3835 = ~( N3712 | N3768 );
	assign N3837 = ~( N3612 | N3768 );
	assign N3899 = ~( N3835 | N3836 );
	assign N4183 = ~( N4058 | N4118 );
	assign N4185 = ~( N3955 | N4118 );
	assign N4245 = ~( N4183 | N4184 );
	assign N4534 = ~( N4411 | N4470 );
	assign N4536 = ~( N4302 | N4470 );
	assign N4595 = ~( N4534 | N4535 );
	assign N4889 = ~( N4766 | N4825 );
	assign N4891 = ~( N4654 | N4825 );
	assign N4950 = ~( N4889 | N4890 );
	assign N5249 = ~( N5124 | N5184 );
	assign N5251 = ~( N5013 | N5184 );
	assign N5312 = ~( N5249 | N5250 );
	assign N5616 = ~( N5486 | N5548 );
	assign N5618 = ~( N5374 | N5548 );
	assign N5676 = ~( N5616 | N5617 );
	assign N5890 = ~( N5789 | N5840 );
	assign N5892 = ~( N5679 | N5840 );
	assign N5938 = ~( N5890 | N5891 );
	assign N6068 = ~( N6011 | N6040 );
	assign N6070 = ~( N5941 | N6040 );
	assign N6094 = ~( N6068 | N6069 );
	assign N1521 = ~( N1323 | N1458 );
	assign N1588 = ~( N1521 | N1522 );
	assign N1839 = ~( N1726 | N1775 );
	assign N1841 = ~( N1640 | N1775 );
	assign N1908 = ~( N1839 | N1840 );
	assign N2164 = ~( N2046 | N2097 );
	assign N2166 = ~( N1959 | N2097 );
	assign N2230 = ~( N2164 | N2165 );
	assign N2491 = ~( N2371 | N2426 );
	assign N2493 = ~( N2281 | N2426 );
	assign N2555 = ~( N2491 | N2492 );
	assign N2821 = ~( N2703 | N2757 );
	assign N2823 = ~( N2607 | N2757 );
	assign N2884 = ~( N2821 | N2822 );
	assign N3155 = ~( N3037 | N3091 );
	assign N3157 = ~( N2938 | N3091 );
	assign N3218 = ~( N3155 | N3156 );
	assign N3494 = ~( N3374 | N3429 );
	assign N3496 = ~( N3276 | N3429 );
	assign N3559 = ~( N3494 | N3495 );
	assign N3840 = ~( N3715 | N3772 );
	assign N3842 = ~( N3616 | N3772 );
	assign N3902 = ~( N3840 | N3841 );
	assign N4188 = ~( N4061 | N4122 );
	assign N4190 = ~( N3959 | N4122 );
	assign N4248 = ~( N4188 | N4189 );
	assign N4539 = ~( N4414 | N4474 );
	assign N4541 = ~( N4306 | N4474 );
	assign N4598 = ~( N4539 | N4540 );
	assign N4894 = ~( N4769 | N4829 );
	assign N4896 = ~( N4658 | N4829 );
	assign N4953 = ~( N4894 | N4895 );
	assign N5254 = ~( N5127 | N5188 );
	assign N5256 = ~( N5017 | N5188 );
	assign N5315 = ~( N5254 | N5255 );
	assign N5552 = ~( N5431 | N5489 );
	assign N5554 = ~( N5318 | N5489 );
	assign N5621 = ~( N5552 | N5553 );
	assign N5844 = ~( N5740 | N5792 );
	assign N5846 = ~( N5624 | N5792 );
	assign N5895 = ~( N5844 | N5845 );
	assign N6044 = ~( N5981 | N6014 );
	assign N6046 = ~( N5898 | N6014 );
	assign N6073 = ~( N6044 | N6045 );
	assign N1526 = ~( N1327 | N1462 );
	assign N1591 = ~( N1526 | N1527 );
	assign N1844 = ~( N1729 | N1779 );
	assign N1846 = ~( N1644 | N1779 );
	assign N1911 = ~( N1844 | N1845 );
	assign N2169 = ~( N2049 | N2101 );
	assign N2171 = ~( N1963 | N2101 );
	assign N2233 = ~( N2169 | N2170 );
	assign N2496 = ~( N2374 | N2430 );
	assign N2498 = ~( N2285 | N2430 );
	assign N2558 = ~( N2496 | N2497 );
	assign N2826 = ~( N2706 | N2761 );
	assign N2828 = ~( N2611 | N2761 );
	assign N2887 = ~( N2826 | N2827 );
	assign N3160 = ~( N3040 | N3095 );
	assign N3162 = ~( N2942 | N3095 );
	assign N3221 = ~( N3160 | N3161 );
	assign N3499 = ~( N3377 | N3433 );
	assign N3501 = ~( N3280 | N3433 );
	assign N3562 = ~( N3499 | N3500 );
	assign N3845 = ~( N3718 | N3776 );
	assign N3847 = ~( N3620 | N3776 );
	assign N3905 = ~( N3845 | N3846 );
	assign N4193 = ~( N4064 | N4126 );
	assign N4195 = ~( N3963 | N4126 );
	assign N4251 = ~( N4193 | N4194 );
	assign N4544 = ~( N4417 | N4478 );
	assign N4546 = ~( N4310 | N4478 );
	assign N4601 = ~( N4544 | N4545 );
	assign N4899 = ~( N4772 | N4833 );
	assign N4901 = ~( N4662 | N4833 );
	assign N4956 = ~( N4899 | N4900 );
	assign N5192 = ~( N5073 | N5130 );
	assign N5194 = ~( N4959 | N5130 );
	assign N5259 = ~( N5192 | N5193 );
	assign N5493 = ~( N5380 | N5434 );
	assign N5495 = ~( N5262 | N5434 );
	assign N5557 = ~( N5493 | N5494 );
	assign N5796 = ~( N5685 | N5743 );
	assign N5798 = ~( N5560 | N5743 );
	assign N5849 = ~( N5796 | N5797 );
	assign N6018 = ~( N5947 | N5984 );
	assign N6020 = ~( N5852 | N5984 );
	assign N6049 = ~( N6018 | N6019 );
	assign N1531 = ~( N1331 | N1466 );
	assign N1594 = ~( N1531 | N1532 );
	assign N1849 = ~( N1732 | N1783 );
	assign N1851 = ~( N1648 | N1783 );
	assign N1914 = ~( N1849 | N1850 );
	assign N2174 = ~( N2052 | N2105 );
	assign N2176 = ~( N1967 | N2105 );
	assign N2236 = ~( N2174 | N2175 );
	assign N2501 = ~( N2377 | N2434 );
	assign N2503 = ~( N2289 | N2434 );
	assign N2561 = ~( N2501 | N2502 );
	assign N2831 = ~( N2709 | N2765 );
	assign N2833 = ~( N2615 | N2765 );
	assign N2890 = ~( N2831 | N2832 );
	assign N3165 = ~( N3043 | N3099 );
	assign N3167 = ~( N2946 | N3099 );
	assign N3224 = ~( N3165 | N3166 );
	assign N3504 = ~( N3380 | N3437 );
	assign N3506 = ~( N3284 | N3437 );
	assign N3565 = ~( N3504 | N3505 );
	assign N3850 = ~( N3721 | N3780 );
	assign N3852 = ~( N3624 | N3780 );
	assign N3908 = ~( N3850 | N3851 );
	assign N4198 = ~( N4067 | N4130 );
	assign N4200 = ~( N3967 | N4130 );
	assign N4254 = ~( N4198 | N4199 );
	assign N4549 = ~( N4420 | N4482 );
	assign N4551 = ~( N4314 | N4482 );
	assign N4604 = ~( N4549 | N4550 );
	assign N4837 = ~( N4718 | N4775 );
	assign N4839 = ~( N4607 | N4775 );
	assign N4904 = ~( N4837 | N4838 );
	assign N5134 = ~( N5023 | N5076 );
	assign N5136 = ~( N4907 | N5076 );
	assign N5197 = ~( N5134 | N5135 );
	assign N5438 = ~( N5324 | N5383 );
	assign N5440 = ~( N5200 | N5383 );
	assign N5498 = ~( N5438 | N5439 );
	assign N5747 = ~( N5630 | N5688 );
	assign N5749 = ~( N5501 | N5688 );
	assign N5801 = ~( N5747 | N5748 );
	assign N5988 = ~( N5904 | N5950 );
	assign N5990 = ~( N5804 | N5950 );
	assign N6023 = ~( N5988 | N5989 );
	assign N1536 = ~( N1335 | N1470 );
	assign N1597 = ~( N1536 | N1537 );
	assign N1854 = ~( N1735 | N1787 );
	assign N1856 = ~( N1652 | N1787 );
	assign N1917 = ~( N1854 | N1855 );
	assign N2179 = ~( N2055 | N2109 );
	assign N2181 = ~( N1971 | N2109 );
	assign N2239 = ~( N2179 | N2180 );
	assign N2506 = ~( N2380 | N2438 );
	assign N2508 = ~( N2293 | N2438 );
	assign N2564 = ~( N2506 | N2507 );
	assign N2836 = ~( N2712 | N2769 );
	assign N2838 = ~( N2619 | N2769 );
	assign N2893 = ~( N2836 | N2837 );
	assign N3170 = ~( N3046 | N3103 );
	assign N3172 = ~( N2950 | N3103 );
	assign N3227 = ~( N3170 | N3171 );
	assign N3509 = ~( N3383 | N3441 );
	assign N3511 = ~( N3288 | N3441 );
	assign N3568 = ~( N3509 | N3510 );
	assign N3855 = ~( N3724 | N3784 );
	assign N3857 = ~( N3628 | N3784 );
	assign N3911 = ~( N3855 | N3856 );
	assign N4203 = ~( N4070 | N4134 );
	assign N4205 = ~( N3971 | N4134 );
	assign N4257 = ~( N4203 | N4204 );
	assign N4486 = ~( N4365 | N4423 );
	assign N4488 = ~( N4260 | N4423 );
	assign N4554 = ~( N4486 | N4487 );
	assign N4779 = ~( N4668 | N4721 );
	assign N4781 = ~( N4557 | N4721 );
	assign N4842 = ~( N4779 | N4780 );
	assign N5080 = ~( N4965 | N5026 );
	assign N5082 = ~( N4845 | N5026 );
	assign N5139 = ~( N5080 | N5081 );
	assign N5387 = ~( N5268 | N5327 );
	assign N5389 = ~( N5142 | N5327 );
	assign N5443 = ~( N5387 | N5388 );
	assign N5692 = ~( N5566 | N5633 );
	assign N5694 = ~( N5446 | N5633 );
	assign N5752 = ~( N5692 | N5693 );
	assign N5954 = ~( N5858 | N5907 );
	assign N5956 = ~( N5755 | N5907 );
	assign N5993 = ~( N5954 | N5955 );
	assign N1541 = ~( N1339 | N1474 );
	assign N1600 = ~( N1541 | N1542 );
	assign N1859 = ~( N1738 | N1791 );
	assign N1861 = ~( N1656 | N1791 );
	assign N1920 = ~( N1859 | N1860 );
	assign N2184 = ~( N2058 | N2113 );
	assign N2186 = ~( N1975 | N2113 );
	assign N2242 = ~( N2184 | N2185 );
	assign N2511 = ~( N2383 | N2442 );
	assign N2513 = ~( N2297 | N2442 );
	assign N2567 = ~( N2511 | N2512 );
	assign N2841 = ~( N2715 | N2773 );
	assign N2843 = ~( N2623 | N2773 );
	assign N2896 = ~( N2841 | N2842 );
	assign N3175 = ~( N3049 | N3107 );
	assign N3177 = ~( N2954 | N3107 );
	assign N3230 = ~( N3175 | N3176 );
	assign N3514 = ~( N3386 | N3445 );
	assign N3516 = ~( N3292 | N3445 );
	assign N3571 = ~( N3514 | N3515 );
	assign N3860 = ~( N3727 | N3788 );
	assign N3862 = ~( N3632 | N3788 );
	assign N3914 = ~( N3860 | N3861 );
	assign N4138 = ~( N4019 | N4073 );
	assign N4140 = ~( N3917 | N4073 );
	assign N4208 = ~( N4138 | N4139 );
	assign N4427 = ~( N4320 | N4368 );
	assign N4429 = ~( N4211 | N4368 );
	assign N4491 = ~( N4427 | N4428 );
	assign N4725 = ~( N4613 | N4671 );
	assign N4727 = ~( N4494 | N4671 );
	assign N4784 = ~( N4725 | N4726 );
	assign N5030 = ~( N4913 | N4968 );
	assign N5032 = ~( N4787 | N4968 );
	assign N5085 = ~( N5030 | N5031 );
	assign N5331 = ~( N5206 | N5271 );
	assign N5333 = ~( N5088 | N5271 );
	assign N5392 = ~( N5331 | N5332 );
	assign N5637 = ~( N5507 | N5569 );
	assign N5639 = ~( N5395 | N5569 );
	assign N5697 = ~( N5637 | N5638 );
	assign N5911 = ~( N5810 | N5861 );
	assign N5913 = ~( N5700 | N5861 );
	assign N5959 = ~( N5911 | N5912 );
	assign N1546 = ~( N1343 | N1478 );
	assign N1603 = ~( N1546 | N1547 );
	assign N1864 = ~( N1741 | N1795 );
	assign N1866 = ~( N1660 | N1795 );
	assign N1923 = ~( N1864 | N1865 );
	assign N2189 = ~( N2061 | N2117 );
	assign N2191 = ~( N1979 | N2117 );
	assign N2245 = ~( N2189 | N2190 );
	assign N2516 = ~( N2386 | N2446 );
	assign N2518 = ~( N2301 | N2446 );
	assign N2570 = ~( N2516 | N2517 );
	assign N2846 = ~( N2718 | N2777 );
	assign N2848 = ~( N2627 | N2777 );
	assign N2899 = ~( N2846 | N2847 );
	assign N3180 = ~( N3052 | N3111 );
	assign N3182 = ~( N2958 | N3111 );
	assign N3233 = ~( N3180 | N3181 );
	assign N3519 = ~( N3389 | N3449 );
	assign N3521 = ~( N3296 | N3449 );
	assign N3574 = ~( N3519 | N3520 );
	assign N3792 = ~( N3678 | N3730 );
	assign N3794 = ~( N3577 | N3730 );
	assign N3865 = ~( N3792 | N3793 );
	assign N4077 = ~( N3977 | N4022 );
	assign N4079 = ~( N3868 | N4022 );
	assign N4143 = ~( N4077 | N4078 );
	assign N4372 = ~( N4266 | N4323 );
	assign N4374 = ~( N4146 | N4323 );
	assign N4432 = ~( N4372 | N4373 );
	assign N4675 = ~( N4563 | N4616 );
	assign N4677 = ~( N4435 | N4616 );
	assign N4730 = ~( N4675 | N4676 );
	assign N4972 = ~( N4851 | N4916 );
	assign N4974 = ~( N4733 | N4916 );
	assign N5035 = ~( N4972 | N4973 );
	assign N5275 = ~( N5148 | N5209 );
	assign N5277 = ~( N5038 | N5209 );
	assign N5336 = ~( N5275 | N5276 );
	assign N5573 = ~( N5452 | N5510 );
	assign N5575 = ~( N5339 | N5510 );
	assign N5642 = ~( N5573 | N5574 );
	assign N5865 = ~( N5761 | N5813 );
	assign N5867 = ~( N5645 | N5813 );
	assign N5916 = ~( N5865 | N5866 );
	assign N1551 = ~( N1347 | N1482 );
	assign N1606 = ~( N1551 | N1552 );
	assign N1869 = ~( N1744 | N1799 );
	assign N1871 = ~( N1664 | N1799 );
	assign N1926 = ~( N1869 | N1870 );
	assign N2194 = ~( N2064 | N2121 );
	assign N2196 = ~( N1983 | N2121 );
	assign N2248 = ~( N2194 | N2195 );
	assign N2521 = ~( N2389 | N2450 );
	assign N2523 = ~( N2305 | N2450 );
	assign N2573 = ~( N2521 | N2522 );
	assign N2851 = ~( N2721 | N2781 );
	assign N2853 = ~( N2631 | N2781 );
	assign N2902 = ~( N2851 | N2852 );
	assign N3185 = ~( N3055 | N3115 );
	assign N3187 = ~( N2962 | N3115 );
	assign N3236 = ~( N3185 | N3186 );
	assign N3453 = ~( N3341 | N3392 );
	assign N3455 = ~( N3239 | N3392 );
	assign N3524 = ~( N3453 | N3454 );
	assign N3734 = ~( N3638 | N3681 );
	assign N3736 = ~( N3527 | N3681 );
	assign N3797 = ~( N3734 | N3735 );
	assign N4026 = ~( N3923 | N3980 );
	assign N4028 = ~( N3800 | N3980 );
	assign N4082 = ~( N4026 | N4027 );
	assign N4327 = ~( N4217 | N4269 );
	assign N4329 = ~( N4085 | N4269 );
	assign N4377 = ~( N4327 | N4328 );
	assign N4620 = ~( N4500 | N4566 );
	assign N4622 = ~( N4380 | N4566 );
	assign N4680 = ~( N4620 | N4621 );
	assign N4920 = ~( N4793 | N4854 );
	assign N4922 = ~( N4683 | N4854 );
	assign N4977 = ~( N4920 | N4921 );
	assign N5213 = ~( N5094 | N5151 );
	assign N5215 = ~( N4980 | N5151 );
	assign N5280 = ~( N5213 | N5214 );
	assign N5514 = ~( N5401 | N5455 );
	assign N5516 = ~( N5283 | N5455 );
	assign N5578 = ~( N5514 | N5515 );
	assign N5817 = ~( N5706 | N5764 );
	assign N5819 = ~( N5581 | N5764 );
	assign N5870 = ~( N5817 | N5818 );
	assign N1556 = ~( N1351 | N1486 );
	assign N1609 = ~( N1556 | N1557 );
	assign N1874 = ~( N1747 | N1803 );
	assign N1876 = ~( N1668 | N1803 );
	assign N1929 = ~( N1874 | N1875 );
	assign N2199 = ~( N2067 | N2125 );
	assign N2201 = ~( N1987 | N2125 );
	assign N2251 = ~( N2199 | N2200 );
	assign N2526 = ~( N2392 | N2454 );
	assign N2528 = ~( N2309 | N2454 );
	assign N2576 = ~( N2526 | N2527 );
	assign N2856 = ~( N2724 | N2785 );
	assign N2858 = ~( N2635 | N2785 );
	assign N2905 = ~( N2856 | N2857 );
	assign N3119 = ~( N3007 | N3058 );
	assign N3121 = ~( N2908 | N3058 );
	assign N3190 = ~( N3119 | N3120 );
	assign N3396 = ~( N3302 | N3344 );
	assign N3398 = ~( N3193 | N3344 );
	assign N3458 = ~( N3396 | N3397 );
	assign N3685 = ~( N3583 | N3641 );
	assign N3687 = ~( N3461 | N3641 );
	assign N3739 = ~( N3685 | N3686 );
	assign N3984 = ~( N3874 | N3926 );
	assign N3986 = ~( N3742 | N3926 );
	assign N4031 = ~( N3984 | N3985 );
	assign N4273 = ~( N4152 | N4220 );
	assign N4275 = ~( N4034 | N4220 );
	assign N4332 = ~( N4273 | N4274 );
	assign N4570 = ~( N4441 | N4503 );
	assign N4572 = ~( N4335 | N4503 );
	assign N4625 = ~( N4570 | N4571 );
	assign N4858 = ~( N4739 | N4796 );
	assign N4860 = ~( N4628 | N4796 );
	assign N4925 = ~( N4858 | N4859 );
	assign N5155 = ~( N5044 | N5097 );
	assign N5157 = ~( N4928 | N5097 );
	assign N5218 = ~( N5155 | N5156 );
	assign N5459 = ~( N5345 | N5404 );
	assign N5461 = ~( N5221 | N5404 );
	assign N5519 = ~( N5459 | N5460 );
	assign N5768 = ~( N5651 | N5709 );
	assign N5770 = ~( N5522 | N5709 );
	assign N5822 = ~( N5768 | N5769 );
	assign N1561 = ~( N1355 | N1490 );
	assign N1612 = ~( N1561 | N1562 );
	assign N1879 = ~( N1750 | N1807 );
	assign N1881 = ~( N1672 | N1807 );
	assign N1932 = ~( N1879 | N1880 );
	assign N2204 = ~( N2070 | N2129 );
	assign N2206 = ~( N1991 | N2129 );
	assign N2254 = ~( N2204 | N2205 );
	assign N2531 = ~( N2395 | N2458 );
	assign N2533 = ~( N2313 | N2458 );
	assign N2579 = ~( N2531 | N2532 );
	assign N2789 = ~( N2675 | N2727 );
	assign N2791 = ~( N2582 | N2727 );
	assign N2861 = ~( N2789 | N2790 );
	assign N3062 = ~( N2968 | N3010 );
	assign N3064 = ~( N2864 | N3010 );
	assign N3124 = ~( N3062 | N3063 );
	assign N3348 = ~( N3245 | N3305 );
	assign N3350 = ~( N3127 | N3305 );
	assign N3401 = ~( N3348 | N3349 );
	assign N3645 = ~( N3533 | N3586 );
	assign N3647 = ~( N3404 | N3586 );
	assign N3690 = ~( N3645 | N3646 );
	assign N3930 = ~( N3806 | N3877 );
	assign N3932 = ~( N3693 | N3877 );
	assign N3989 = ~( N3930 | N3931 );
	assign N4224 = ~( N4091 | N4155 );
	assign N4226 = ~( N3992 | N4155 );
	assign N4278 = ~( N4224 | N4225 );
	assign N4507 = ~( N4386 | N4444 );
	assign N4509 = ~( N4281 | N4444 );
	assign N4575 = ~( N4507 | N4508 );
	assign N4800 = ~( N4689 | N4742 );
	assign N4802 = ~( N4578 | N4742 );
	assign N4863 = ~( N4800 | N4801 );
	assign N5101 = ~( N4986 | N5047 );
	assign N5103 = ~( N4866 | N5047 );
	assign N5160 = ~( N5101 | N5102 );
	assign N5408 = ~( N5289 | N5348 );
	assign N5410 = ~( N5163 | N5348 );
	assign N5464 = ~( N5408 | N5409 );
	assign N5713 = ~( N5587 | N5654 );
	assign N5715 = ~( N5467 | N5654 );
	assign N5773 = ~( N5713 | N5714 );
	assign N1566 = ~( N1359 | N1494 );
	assign N1615 = ~( N1566 | N1567 );
	assign N1884 = ~( N1753 | N1811 );
	assign N1886 = ~( N1676 | N1811 );
	assign N1935 = ~( N1884 | N1885 );
	assign N2209 = ~( N2073 | N2133 );
	assign N2211 = ~( N1995 | N2133 );
	assign N2257 = ~( N2209 | N2210 );
	assign N2462 = ~( N2350 | N2398 );
	assign N2464 = ~( N2260 | N2398 );
	assign N2536 = ~( N2462 | N2463 );
	assign N2731 = ~( N2641 | N2678 );
	assign N2733 = ~( N2539 | N2678 );
	assign N2794 = ~( N2731 | N2732 );
	assign N3014 = ~( N2914 | N2971 );
	assign N3016 = ~( N2797 | N2971 );
	assign N3067 = ~( N3014 | N3015 );
	assign N3309 = ~( N3199 | N3248 );
	assign N3311 = ~( N3070 | N3248 );
	assign N3353 = ~( N3309 | N3310 );
	assign N3590 = ~( N3467 | N3536 );
	assign N3592 = ~( N3356 | N3536 );
	assign N3650 = ~( N3590 | N3591 );
	assign N3881 = ~( N3748 | N3809 );
	assign N3883 = ~( N3653 | N3809 );
	assign N3935 = ~( N3881 | N3882 );
	assign N4159 = ~( N4040 | N4094 );
	assign N4161 = ~( N3938 | N4094 );
	assign N4229 = ~( N4159 | N4160 );
	assign N4448 = ~( N4341 | N4389 );
	assign N4450 = ~( N4232 | N4389 );
	assign N4512 = ~( N4448 | N4449 );
	assign N4746 = ~( N4634 | N4692 );
	assign N4748 = ~( N4515 | N4692 );
	assign N4805 = ~( N4746 | N4747 );
	assign N5051 = ~( N4934 | N4989 );
	assign N5053 = ~( N4808 | N4989 );
	assign N5106 = ~( N5051 | N5052 );
	assign N5352 = ~( N5227 | N5292 );
	assign N5354 = ~( N5109 | N5292 );
	assign N5413 = ~( N5352 | N5353 );
	assign N5658 = ~( N5528 | N5590 );
	assign N5660 = ~( N5416 | N5590 );
	assign N5718 = ~( N5658 | N5659 );
	assign N1571 = ~( N1363 | N1498 );
	assign N1618 = ~( N1571 | N1572 );
	assign N1889 = ~( N1756 | N1815 );
	assign N1891 = ~( N1680 | N1815 );
	assign N1938 = ~( N1889 | N1890 );
	assign N2137 = ~( N2030 | N2076 );
	assign N2139 = ~( N1941 | N2076 );
	assign N2214 = ~( N2137 | N2138 );
	assign N2402 = ~( N2319 | N2353 );
	assign N2404 = ~( N2217 | N2353 );
	assign N2467 = ~( N2402 | N2403 );
	assign N2682 = ~( N2588 | N2644 );
	assign N2684 = ~( N2470 | N2644 );
	assign N2736 = ~( N2682 | N2683 );
	assign N2975 = ~( N2870 | N2917 );
	assign N2977 = ~( N2739 | N2917 );
	assign N3019 = ~( N2975 | N2976 );
	assign N3252 = ~( N3133 | N3202 );
	assign N3254 = ~( N3022 | N3202 );
	assign N3314 = ~( N3252 | N3253 );
	assign N3540 = ~( N3410 | N3470 );
	assign N3542 = ~( N3317 | N3470 );
	assign N3595 = ~( N3540 | N3541 );
	assign N3813 = ~( N3699 | N3751 );
	assign N3815 = ~( N3598 | N3751 );
	assign N3886 = ~( N3813 | N3814 );
	assign N4098 = ~( N3998 | N4043 );
	assign N4100 = ~( N3889 | N4043 );
	assign N4164 = ~( N4098 | N4099 );
	assign N4393 = ~( N4287 | N4344 );
	assign N4395 = ~( N4167 | N4344 );
	assign N4453 = ~( N4393 | N4394 );
	assign N4696 = ~( N4584 | N4637 );
	assign N4698 = ~( N4456 | N4637 );
	assign N4751 = ~( N4696 | N4697 );
	assign N4993 = ~( N4872 | N4937 );
	assign N4995 = ~( N4754 | N4937 );
	assign N5056 = ~( N4993 | N4994 );
	assign N5296 = ~( N5169 | N5230 );
	assign N5298 = ~( N5059 | N5230 );
	assign N5357 = ~( N5296 | N5297 );
	assign N5594 = ~( N5473 | N5531 );
	assign N5596 = ~( N5360 | N5531 );
	assign N5663 = ~( N5594 | N5595 );
	assign N1576 = ~( N1367 | N1502 );
	assign N1621 = ~( N1576 | N1577 );
	assign N1819 = ~( N1714 | N1759 );
	assign N1821 = ~( N1624 | N1759 );
	assign N1894 = ~( N1819 | N1820 );
	assign N2080 = ~( N2001 | N2033 );
	assign N2082 = ~( N1897 | N2033 );
	assign N2142 = ~( N2080 | N2081 );
	assign N2357 = ~( N2266 | N2322 );
	assign N2359 = ~( N2145 | N2322 );
	assign N2407 = ~( N2357 | N2358 );
	assign N2648 = ~( N2545 | N2591 );
	assign N2650 = ~( N2410 | N2591 );
	assign N2687 = ~( N2648 | N2649 );
	assign N2921 = ~( N2803 | N2873 );
	assign N2923 = ~( N2690 | N2873 );
	assign N2980 = ~( N2921 | N2922 );
	assign N3206 = ~( N3076 | N3136 );
	assign N3208 = ~( N2983 | N3136 );
	assign N3257 = ~( N3206 | N3207 );
	assign N3474 = ~( N3362 | N3413 );
	assign N3476 = ~( N3260 | N3413 );
	assign N3545 = ~( N3474 | N3475 );
	assign N3755 = ~( N3659 | N3702 );
	assign N3757 = ~( N3548 | N3702 );
	assign N3818 = ~( N3755 | N3756 );
	assign N4047 = ~( N3944 | N4001 );
	assign N4049 = ~( N3821 | N4001 );
	assign N4103 = ~( N4047 | N4048 );
	assign N4348 = ~( N4238 | N4290 );
	assign N4350 = ~( N4106 | N4290 );
	assign N4398 = ~( N4348 | N4349 );
	assign N4641 = ~( N4521 | N4587 );
	assign N4643 = ~( N4401 | N4587 );
	assign N4701 = ~( N4641 | N4642 );
	assign N4941 = ~( N4814 | N4875 );
	assign N4943 = ~( N4704 | N4875 );
	assign N4998 = ~( N4941 | N4942 );
	assign N5234 = ~( N5115 | N5172 );
	assign N5236 = ~( N5001 | N5172 );
	assign N5301 = ~( N5234 | N5235 );
	assign N5535 = ~( N5422 | N5476 );
	assign N5537 = ~( N5304 | N5476 );
	assign N5599 = ~( N5535 | N5536 );
	assign N1685 = ~( N1624 | N1576 );
	assign N1714 = ~( N1684 | N1685 );
	assign N1946 = ~( N1897 | N1821 );
	assign N2001 = ~( N1945 | N1946 );
	assign N2222 = ~( N2145 | N2082 );
	assign N2266 = ~( N2221 | N2222 );
	assign N2475 = ~( N2410 | N2359 );
	assign N2545 = ~( N2474 | N2475 );
	assign N2744 = ~( N2690 | N2650 );
	assign N2803 = ~( N2743 | N2744 );
	assign N3027 = ~( N2983 | N2923 );
	assign N3076 = ~( N3026 | N3027 );
	assign N3322 = ~( N3260 | N3208 );
	assign N3362 = ~( N3321 | N3322 );
	assign N3603 = ~( N3548 | N3476 );
	assign N3659 = ~( N3602 | N3603 );
	assign N3894 = ~( N3821 | N3757 );
	assign N3944 = ~( N3893 | N3894 );
	assign N4172 = ~( N4106 | N4049 );
	assign N4238 = ~( N4171 | N4172 );
	assign N4461 = ~( N4401 | N4350 );
	assign N4521 = ~( N4460 | N4461 );
	assign N4759 = ~( N4704 | N4643 );
	assign N4814 = ~( N4758 | N4759 );
	assign N5064 = ~( N5001 | N4943 );
	assign N5115 = ~( N5063 | N5064 );
	assign N5365 = ~( N5304 | N5236 );
	assign N5422 = ~( N5364 | N5365 );
	assign N5671 = ~( N5602 | N5537 );
	assign N6287 = ~( N5602 | N6281 );
	assign N5727 = ~( N5670 | N5671 );
	assign N1628 = ~( N1582 | N1506 );
	assign N1687 = ~( N1628 | N1506 );
	assign N1947 = ~( N1902 | N1826 );
	assign N2005 = ~( N1947 | N1826 );
	assign N2269 = ~( N2224 | N2151 );
	assign N2327 = ~( N2269 | N2151 );
	assign N2595 = ~( N2549 | N2478 );
	assign N2654 = ~( N2595 | N2478 );
	assign N2926 = ~( N2878 | N2808 );
	assign N2988 = ~( N2926 | N2808 );
	assign N3264 = ~( N3212 | N3142 );
	assign N3324 = ~( N3264 | N3142 );
	assign N3604 = ~( N3553 | N3481 );
	assign N3663 = ~( N3604 | N3481 );
	assign N3947 = ~( N3896 | N3827 );
	assign N4006 = ~( N3947 | N3827 );
	assign N4294 = ~( N4242 | N4175 );
	assign N4354 = ~( N4294 | N4175 );
	assign N4646 = ~( N4592 | N4526 );
	assign N4709 = ~( N4646 | N4526 );
	assign N5005 = ~( N4947 | N4881 );
	assign N5066 = ~( N5005 | N4881 );
	assign N5366 = ~( N5309 | N5241 );
	assign N5426 = ~( N5366 | N5241 );
	assign N5730 = ~( N5673 | N5608 );
	assign N5786 = ~( N5730 | N5608 );
	assign N6005 = ~( N5972 | N5930 );
	assign N6036 = ~( N6005 | N5930 );
	assign N6124 = ~( N6111 | N6108 );
	assign N6134 = ~( N6124 | N6108 );
	assign N1632 = ~( N1585 | N1511 );
	assign N1689 = ~( N1632 | N1511 );
	assign N1686 = ~( N1582 | N1628 );
	assign N1951 = ~( N1905 | N1831 );
	assign N2007 = ~( N1951 | N1831 );
	assign N2004 = ~( N1902 | N1947 );
	assign N2273 = ~( N2227 | N2156 );
	assign N2329 = ~( N2273 | N2156 );
	assign N2326 = ~( N2224 | N2269 );
	assign N2599 = ~( N2552 | N2483 );
	assign N2656 = ~( N2599 | N2483 );
	assign N2653 = ~( N2549 | N2595 );
	assign N2930 = ~( N2881 | N2813 );
	assign N2990 = ~( N2930 | N2813 );
	assign N2987 = ~( N2878 | N2926 );
	assign N3268 = ~( N3215 | N3147 );
	assign N3326 = ~( N3268 | N3147 );
	assign N3323 = ~( N3212 | N3264 );
	assign N3608 = ~( N3556 | N3486 );
	assign N3665 = ~( N3608 | N3486 );
	assign N3662 = ~( N3553 | N3604 );
	assign N3951 = ~( N3899 | N3832 );
	assign N4008 = ~( N3951 | N3832 );
	assign N4005 = ~( N3896 | N3947 );
	assign N4298 = ~( N4245 | N4180 );
	assign N4356 = ~( N4298 | N4180 );
	assign N4353 = ~( N4242 | N4294 );
	assign N4650 = ~( N4595 | N4531 );
	assign N4711 = ~( N4650 | N4531 );
	assign N4708 = ~( N4592 | N4646 );
	assign N5009 = ~( N4950 | N4886 );
	assign N5068 = ~( N5009 | N4886 );
	assign N5065 = ~( N4947 | N5005 );
	assign N5370 = ~( N5312 | N5246 );
	assign N5428 = ~( N5370 | N5246 );
	assign N5425 = ~( N5309 | N5366 );
	assign N5734 = ~( N5676 | N5613 );
	assign N5788 = ~( N5734 | N5613 );
	assign N5785 = ~( N5673 | N5730 );
	assign N5975 = ~( N5938 | N5935 );
	assign N6010 = ~( N5975 | N5935 );
	assign N6035 = ~( N5972 | N6005 );
	assign N6114 = ~( N6094 | N6091 );
	assign N6129 = ~( N6114 | N6091 );
	assign N6133 = ~( N6111 | N6124 );
	assign N1636 = ~( N1588 | N1516 );
	assign N1691 = ~( N1636 | N1516 );
	assign N1688 = ~( N1585 | N1632 );
	assign N1955 = ~( N1908 | N1836 );
	assign N2009 = ~( N1955 | N1836 );
	assign N2006 = ~( N1905 | N1951 );
	assign N2277 = ~( N2230 | N2161 );
	assign N2331 = ~( N2277 | N2161 );
	assign N2328 = ~( N2227 | N2273 );
	assign N2603 = ~( N2555 | N2488 );
	assign N2658 = ~( N2603 | N2488 );
	assign N2655 = ~( N2552 | N2599 );
	assign N2934 = ~( N2884 | N2818 );
	assign N2992 = ~( N2934 | N2818 );
	assign N2989 = ~( N2881 | N2930 );
	assign N3272 = ~( N3218 | N3152 );
	assign N3328 = ~( N3272 | N3152 );
	assign N3325 = ~( N3215 | N3268 );
	assign N3612 = ~( N3559 | N3491 );
	assign N3667 = ~( N3612 | N3491 );
	assign N3664 = ~( N3556 | N3608 );
	assign N3955 = ~( N3902 | N3837 );
	assign N4010 = ~( N3955 | N3837 );
	assign N4007 = ~( N3899 | N3951 );
	assign N4302 = ~( N4248 | N4185 );
	assign N4358 = ~( N4302 | N4185 );
	assign N4355 = ~( N4245 | N4298 );
	assign N4654 = ~( N4598 | N4536 );
	assign N4713 = ~( N4654 | N4536 );
	assign N4710 = ~( N4595 | N4650 );
	assign N5013 = ~( N4953 | N4891 );
	assign N5070 = ~( N5013 | N4891 );
	assign N5067 = ~( N4950 | N5009 );
	assign N5374 = ~( N5315 | N5251 );
	assign N5430 = ~( N5374 | N5251 );
	assign N5427 = ~( N5312 | N5370 );
	assign N5679 = ~( N5621 | N5618 );
	assign N5739 = ~( N5679 | N5618 );
	assign N5787 = ~( N5676 | N5734 );
	assign N5941 = ~( N5895 | N5892 );
	assign N5980 = ~( N5941 | N5892 );
	assign N6009 = ~( N5938 | N5975 );
	assign N6097 = ~( N6073 | N6070 );
	assign N6119 = ~( N6097 | N6070 );
	assign N6128 = ~( N6094 | N6114 );
	assign N1640 = ~( N1591 | N1521 );
	assign N1693 = ~( N1640 | N1521 );
	assign N1690 = ~( N1588 | N1636 );
	assign N1959 = ~( N1911 | N1841 );
	assign N2011 = ~( N1959 | N1841 );
	assign N2008 = ~( N1908 | N1955 );
	assign N2281 = ~( N2233 | N2166 );
	assign N2333 = ~( N2281 | N2166 );
	assign N2330 = ~( N2230 | N2277 );
	assign N2607 = ~( N2558 | N2493 );
	assign N2660 = ~( N2607 | N2493 );
	assign N2657 = ~( N2555 | N2603 );
	assign N2938 = ~( N2887 | N2823 );
	assign N2994 = ~( N2938 | N2823 );
	assign N2991 = ~( N2884 | N2934 );
	assign N3276 = ~( N3221 | N3157 );
	assign N3330 = ~( N3276 | N3157 );
	assign N3327 = ~( N3218 | N3272 );
	assign N3616 = ~( N3562 | N3496 );
	assign N3669 = ~( N3616 | N3496 );
	assign N3666 = ~( N3559 | N3612 );
	assign N3959 = ~( N3905 | N3842 );
	assign N4012 = ~( N3959 | N3842 );
	assign N4009 = ~( N3902 | N3955 );
	assign N4306 = ~( N4251 | N4190 );
	assign N4360 = ~( N4306 | N4190 );
	assign N4357 = ~( N4248 | N4302 );
	assign N4658 = ~( N4601 | N4541 );
	assign N4715 = ~( N4658 | N4541 );
	assign N4712 = ~( N4598 | N4654 );
	assign N5017 = ~( N4956 | N4896 );
	assign N5072 = ~( N5017 | N4896 );
	assign N5069 = ~( N4953 | N5013 );
	assign N5318 = ~( N5259 | N5256 );
	assign N5379 = ~( N5318 | N5256 );
	assign N5429 = ~( N5315 | N5374 );
	assign N5624 = ~( N5557 | N5554 );
	assign N5684 = ~( N5624 | N5554 );
	assign N5738 = ~( N5621 | N5679 );
	assign N5898 = ~( N5849 | N5846 );
	assign N5946 = ~( N5898 | N5846 );
	assign N5979 = ~( N5895 | N5941 );
	assign N6076 = ~( N6049 | N6046 );
	assign N6102 = ~( N6076 | N6046 );
	assign N6118 = ~( N6073 | N6097 );
	assign N1644 = ~( N1594 | N1526 );
	assign N1695 = ~( N1644 | N1526 );
	assign N1692 = ~( N1591 | N1640 );
	assign N1963 = ~( N1914 | N1846 );
	assign N2013 = ~( N1963 | N1846 );
	assign N2010 = ~( N1911 | N1959 );
	assign N2285 = ~( N2236 | N2171 );
	assign N2335 = ~( N2285 | N2171 );
	assign N2332 = ~( N2233 | N2281 );
	assign N2611 = ~( N2561 | N2498 );
	assign N2662 = ~( N2611 | N2498 );
	assign N2659 = ~( N2558 | N2607 );
	assign N2942 = ~( N2890 | N2828 );
	assign N2996 = ~( N2942 | N2828 );
	assign N2993 = ~( N2887 | N2938 );
	assign N3280 = ~( N3224 | N3162 );
	assign N3332 = ~( N3280 | N3162 );
	assign N3329 = ~( N3221 | N3276 );
	assign N3620 = ~( N3565 | N3501 );
	assign N3671 = ~( N3620 | N3501 );
	assign N3668 = ~( N3562 | N3616 );
	assign N3963 = ~( N3908 | N3847 );
	assign N4014 = ~( N3963 | N3847 );
	assign N4011 = ~( N3905 | N3959 );
	assign N4310 = ~( N4254 | N4195 );
	assign N4362 = ~( N4310 | N4195 );
	assign N4359 = ~( N4251 | N4306 );
	assign N4662 = ~( N4604 | N4546 );
	assign N4717 = ~( N4662 | N4546 );
	assign N4714 = ~( N4601 | N4658 );
	assign N4959 = ~( N4904 | N4901 );
	assign N5022 = ~( N4959 | N4901 );
	assign N5071 = ~( N4956 | N5017 );
	assign N5262 = ~( N5197 | N5194 );
	assign N5323 = ~( N5262 | N5194 );
	assign N5378 = ~( N5259 | N5318 );
	assign N5560 = ~( N5498 | N5495 );
	assign N5629 = ~( N5560 | N5495 );
	assign N5683 = ~( N5557 | N5624 );
	assign N5852 = ~( N5801 | N5798 );
	assign N5903 = ~( N5852 | N5798 );
	assign N5945 = ~( N5849 | N5898 );
	assign N6052 = ~( N6023 | N6020 );
	assign N6081 = ~( N6052 | N6020 );
	assign N6101 = ~( N6049 | N6076 );
	assign N1648 = ~( N1597 | N1531 );
	assign N1697 = ~( N1648 | N1531 );
	assign N1694 = ~( N1594 | N1644 );
	assign N1967 = ~( N1917 | N1851 );
	assign N2015 = ~( N1967 | N1851 );
	assign N2012 = ~( N1914 | N1963 );
	assign N2289 = ~( N2239 | N2176 );
	assign N2337 = ~( N2289 | N2176 );
	assign N2334 = ~( N2236 | N2285 );
	assign N2615 = ~( N2564 | N2503 );
	assign N2664 = ~( N2615 | N2503 );
	assign N2661 = ~( N2561 | N2611 );
	assign N2946 = ~( N2893 | N2833 );
	assign N2998 = ~( N2946 | N2833 );
	assign N2995 = ~( N2890 | N2942 );
	assign N3284 = ~( N3227 | N3167 );
	assign N3334 = ~( N3284 | N3167 );
	assign N3331 = ~( N3224 | N3280 );
	assign N3624 = ~( N3568 | N3506 );
	assign N3673 = ~( N3624 | N3506 );
	assign N3670 = ~( N3565 | N3620 );
	assign N3967 = ~( N3911 | N3852 );
	assign N4016 = ~( N3967 | N3852 );
	assign N4013 = ~( N3908 | N3963 );
	assign N4314 = ~( N4257 | N4200 );
	assign N4364 = ~( N4314 | N4200 );
	assign N4361 = ~( N4254 | N4310 );
	assign N4607 = ~( N4554 | N4551 );
	assign N4667 = ~( N4607 | N4551 );
	assign N4716 = ~( N4604 | N4662 );
	assign N4907 = ~( N4842 | N4839 );
	assign N4964 = ~( N4907 | N4839 );
	assign N5021 = ~( N4904 | N4959 );
	assign N5200 = ~( N5139 | N5136 );
	assign N5267 = ~( N5200 | N5136 );
	assign N5322 = ~( N5197 | N5262 );
	assign N5501 = ~( N5443 | N5440 );
	assign N5565 = ~( N5501 | N5440 );
	assign N5628 = ~( N5498 | N5560 );
	assign N5804 = ~( N5752 | N5749 );
	assign N5857 = ~( N5804 | N5749 );
	assign N5902 = ~( N5801 | N5852 );
	assign N6026 = ~( N5993 | N5990 );
	assign N6057 = ~( N6026 | N5990 );
	assign N6080 = ~( N6023 | N6052 );
	assign N1652 = ~( N1600 | N1536 );
	assign N1699 = ~( N1652 | N1536 );
	assign N1696 = ~( N1597 | N1648 );
	assign N1971 = ~( N1920 | N1856 );
	assign N2017 = ~( N1971 | N1856 );
	assign N2014 = ~( N1917 | N1967 );
	assign N2293 = ~( N2242 | N2181 );
	assign N2339 = ~( N2293 | N2181 );
	assign N2336 = ~( N2239 | N2289 );
	assign N2619 = ~( N2567 | N2508 );
	assign N2666 = ~( N2619 | N2508 );
	assign N2663 = ~( N2564 | N2615 );
	assign N2950 = ~( N2896 | N2838 );
	assign N3000 = ~( N2950 | N2838 );
	assign N2997 = ~( N2893 | N2946 );
	assign N3288 = ~( N3230 | N3172 );
	assign N3336 = ~( N3288 | N3172 );
	assign N3333 = ~( N3227 | N3284 );
	assign N3628 = ~( N3571 | N3511 );
	assign N3675 = ~( N3628 | N3511 );
	assign N3672 = ~( N3568 | N3624 );
	assign N3971 = ~( N3914 | N3857 );
	assign N4018 = ~( N3971 | N3857 );
	assign N4015 = ~( N3911 | N3967 );
	assign N4260 = ~( N4208 | N4205 );
	assign N4319 = ~( N4260 | N4205 );
	assign N4363 = ~( N4257 | N4314 );
	assign N4557 = ~( N4491 | N4488 );
	assign N4612 = ~( N4557 | N4488 );
	assign N4666 = ~( N4554 | N4607 );
	assign N4845 = ~( N4784 | N4781 );
	assign N4912 = ~( N4845 | N4781 );
	assign N4963 = ~( N4842 | N4907 );
	assign N5142 = ~( N5085 | N5082 );
	assign N5205 = ~( N5142 | N5082 );
	assign N5266 = ~( N5139 | N5200 );
	assign N5446 = ~( N5392 | N5389 );
	assign N5506 = ~( N5446 | N5389 );
	assign N5564 = ~( N5443 | N5501 );
	assign N5755 = ~( N5697 | N5694 );
	assign N5809 = ~( N5755 | N5694 );
	assign N5856 = ~( N5752 | N5804 );
	assign N5996 = ~( N5959 | N5956 );
	assign N6031 = ~( N5996 | N5956 );
	assign N6056 = ~( N5993 | N6026 );
	assign N1656 = ~( N1603 | N1541 );
	assign N1701 = ~( N1656 | N1541 );
	assign N1698 = ~( N1600 | N1652 );
	assign N1975 = ~( N1923 | N1861 );
	assign N2019 = ~( N1975 | N1861 );
	assign N2016 = ~( N1920 | N1971 );
	assign N2297 = ~( N2245 | N2186 );
	assign N2341 = ~( N2297 | N2186 );
	assign N2338 = ~( N2242 | N2293 );
	assign N2623 = ~( N2570 | N2513 );
	assign N2668 = ~( N2623 | N2513 );
	assign N2665 = ~( N2567 | N2619 );
	assign N2954 = ~( N2899 | N2843 );
	assign N3002 = ~( N2954 | N2843 );
	assign N2999 = ~( N2896 | N2950 );
	assign N3292 = ~( N3233 | N3177 );
	assign N3338 = ~( N3292 | N3177 );
	assign N3335 = ~( N3230 | N3288 );
	assign N3632 = ~( N3574 | N3516 );
	assign N3677 = ~( N3632 | N3516 );
	assign N3674 = ~( N3571 | N3628 );
	assign N3917 = ~( N3865 | N3862 );
	assign N3976 = ~( N3917 | N3862 );
	assign N4017 = ~( N3914 | N3971 );
	assign N4211 = ~( N4143 | N4140 );
	assign N4265 = ~( N4211 | N4140 );
	assign N4318 = ~( N4208 | N4260 );
	assign N4494 = ~( N4432 | N4429 );
	assign N4562 = ~( N4494 | N4429 );
	assign N4611 = ~( N4491 | N4557 );
	assign N4787 = ~( N4730 | N4727 );
	assign N4850 = ~( N4787 | N4727 );
	assign N4911 = ~( N4784 | N4845 );
	assign N5088 = ~( N5035 | N5032 );
	assign N5147 = ~( N5088 | N5032 );
	assign N5204 = ~( N5085 | N5142 );
	assign N5395 = ~( N5336 | N5333 );
	assign N5451 = ~( N5395 | N5333 );
	assign N5505 = ~( N5392 | N5446 );
	assign N5700 = ~( N5642 | N5639 );
	assign N5760 = ~( N5700 | N5639 );
	assign N5808 = ~( N5697 | N5755 );
	assign N5962 = ~( N5916 | N5913 );
	assign N6001 = ~( N5962 | N5913 );
	assign N6030 = ~( N5959 | N5996 );
	assign N1660 = ~( N1606 | N1546 );
	assign N1703 = ~( N1660 | N1546 );
	assign N1700 = ~( N1603 | N1656 );
	assign N1979 = ~( N1926 | N1866 );
	assign N2021 = ~( N1979 | N1866 );
	assign N2018 = ~( N1923 | N1975 );
	assign N2301 = ~( N2248 | N2191 );
	assign N2343 = ~( N2301 | N2191 );
	assign N2340 = ~( N2245 | N2297 );
	assign N2627 = ~( N2573 | N2518 );
	assign N2670 = ~( N2627 | N2518 );
	assign N2667 = ~( N2570 | N2623 );
	assign N2958 = ~( N2902 | N2848 );
	assign N3004 = ~( N2958 | N2848 );
	assign N3001 = ~( N2899 | N2954 );
	assign N3296 = ~( N3236 | N3182 );
	assign N3340 = ~( N3296 | N3182 );
	assign N3337 = ~( N3233 | N3292 );
	assign N3577 = ~( N3524 | N3521 );
	assign N3637 = ~( N3577 | N3521 );
	assign N3676 = ~( N3574 | N3632 );
	assign N3868 = ~( N3797 | N3794 );
	assign N3922 = ~( N3868 | N3794 );
	assign N3975 = ~( N3865 | N3917 );
	assign N4146 = ~( N4082 | N4079 );
	assign N4216 = ~( N4146 | N4079 );
	assign N4264 = ~( N4143 | N4211 );
	assign N4435 = ~( N4377 | N4374 );
	assign N4499 = ~( N4435 | N4374 );
	assign N4561 = ~( N4432 | N4494 );
	assign N4733 = ~( N4680 | N4677 );
	assign N4792 = ~( N4733 | N4677 );
	assign N4849 = ~( N4730 | N4787 );
	assign N5038 = ~( N4977 | N4974 );
	assign N5093 = ~( N5038 | N4974 );
	assign N5146 = ~( N5035 | N5088 );
	assign N5339 = ~( N5280 | N5277 );
	assign N5400 = ~( N5339 | N5277 );
	assign N5450 = ~( N5336 | N5395 );
	assign N5645 = ~( N5578 | N5575 );
	assign N5705 = ~( N5645 | N5575 );
	assign N5759 = ~( N5642 | N5700 );
	assign N5919 = ~( N5870 | N5867 );
	assign N5967 = ~( N5919 | N5867 );
	assign N6000 = ~( N5916 | N5962 );
	assign N1664 = ~( N1609 | N1551 );
	assign N1705 = ~( N1664 | N1551 );
	assign N1702 = ~( N1606 | N1660 );
	assign N1983 = ~( N1929 | N1871 );
	assign N2023 = ~( N1983 | N1871 );
	assign N2020 = ~( N1926 | N1979 );
	assign N2305 = ~( N2251 | N2196 );
	assign N2345 = ~( N2305 | N2196 );
	assign N2342 = ~( N2248 | N2301 );
	assign N2631 = ~( N2576 | N2523 );
	assign N2672 = ~( N2631 | N2523 );
	assign N2669 = ~( N2573 | N2627 );
	assign N2962 = ~( N2905 | N2853 );
	assign N3006 = ~( N2962 | N2853 );
	assign N3003 = ~( N2902 | N2958 );
	assign N3239 = ~( N3190 | N3187 );
	assign N3301 = ~( N3239 | N3187 );
	assign N3339 = ~( N3236 | N3296 );
	assign N3527 = ~( N3458 | N3455 );
	assign N3582 = ~( N3527 | N3455 );
	assign N3636 = ~( N3524 | N3577 );
	assign N3800 = ~( N3739 | N3736 );
	assign N3873 = ~( N3800 | N3736 );
	assign N3921 = ~( N3797 | N3868 );
	assign N4085 = ~( N4031 | N4028 );
	assign N4151 = ~( N4085 | N4028 );
	assign N4215 = ~( N4082 | N4146 );
	assign N4380 = ~( N4332 | N4329 );
	assign N4440 = ~( N4380 | N4329 );
	assign N4498 = ~( N4377 | N4435 );
	assign N4683 = ~( N4625 | N4622 );
	assign N4738 = ~( N4683 | N4622 );
	assign N4791 = ~( N4680 | N4733 );
	assign N4980 = ~( N4925 | N4922 );
	assign N5043 = ~( N4980 | N4922 );
	assign N5092 = ~( N4977 | N5038 );
	assign N5283 = ~( N5218 | N5215 );
	assign N5344 = ~( N5283 | N5215 );
	assign N5399 = ~( N5280 | N5339 );
	assign N5581 = ~( N5519 | N5516 );
	assign N5650 = ~( N5581 | N5516 );
	assign N5704 = ~( N5578 | N5645 );
	assign N5873 = ~( N5822 | N5819 );
	assign N5924 = ~( N5873 | N5819 );
	assign N5966 = ~( N5870 | N5919 );
	assign N1668 = ~( N1612 | N1556 );
	assign N1707 = ~( N1668 | N1556 );
	assign N1704 = ~( N1609 | N1664 );
	assign N1987 = ~( N1932 | N1876 );
	assign N2025 = ~( N1987 | N1876 );
	assign N2022 = ~( N1929 | N1983 );
	assign N2309 = ~( N2254 | N2201 );
	assign N2347 = ~( N2309 | N2201 );
	assign N2344 = ~( N2251 | N2305 );
	assign N2635 = ~( N2579 | N2528 );
	assign N2674 = ~( N2635 | N2528 );
	assign N2671 = ~( N2576 | N2631 );
	assign N2908 = ~( N2861 | N2858 );
	assign N2967 = ~( N2908 | N2858 );
	assign N3005 = ~( N2905 | N2962 );
	assign N3193 = ~( N3124 | N3121 );
	assign N3244 = ~( N3193 | N3121 );
	assign N3300 = ~( N3190 | N3239 );
	assign N3461 = ~( N3401 | N3398 );
	assign N3532 = ~( N3461 | N3398 );
	assign N3581 = ~( N3458 | N3527 );
	assign N3742 = ~( N3690 | N3687 );
	assign N3805 = ~( N3742 | N3687 );
	assign N3872 = ~( N3739 | N3800 );
	assign N4034 = ~( N3989 | N3986 );
	assign N4090 = ~( N4034 | N3986 );
	assign N4150 = ~( N4031 | N4085 );
	assign N4335 = ~( N4278 | N4275 );
	assign N4385 = ~( N4335 | N4275 );
	assign N4439 = ~( N4332 | N4380 );
	assign N4628 = ~( N4575 | N4572 );
	assign N4688 = ~( N4628 | N4572 );
	assign N4737 = ~( N4625 | N4683 );
	assign N4928 = ~( N4863 | N4860 );
	assign N4985 = ~( N4928 | N4860 );
	assign N5042 = ~( N4925 | N4980 );
	assign N5221 = ~( N5160 | N5157 );
	assign N5288 = ~( N5221 | N5157 );
	assign N5343 = ~( N5218 | N5283 );
	assign N5522 = ~( N5464 | N5461 );
	assign N5586 = ~( N5522 | N5461 );
	assign N5649 = ~( N5519 | N5581 );
	assign N5825 = ~( N5773 | N5770 );
	assign N5878 = ~( N5825 | N5770 );
	assign N5923 = ~( N5822 | N5873 );
	assign N1672 = ~( N1615 | N1561 );
	assign N1709 = ~( N1672 | N1561 );
	assign N1706 = ~( N1612 | N1668 );
	assign N1991 = ~( N1935 | N1881 );
	assign N2027 = ~( N1991 | N1881 );
	assign N2024 = ~( N1932 | N1987 );
	assign N2313 = ~( N2257 | N2206 );
	assign N2349 = ~( N2313 | N2206 );
	assign N2346 = ~( N2254 | N2309 );
	assign N2582 = ~( N2536 | N2533 );
	assign N2640 = ~( N2582 | N2533 );
	assign N2673 = ~( N2579 | N2635 );
	assign N2864 = ~( N2794 | N2791 );
	assign N2913 = ~( N2864 | N2791 );
	assign N2966 = ~( N2861 | N2908 );
	assign N3127 = ~( N3067 | N3064 );
	assign N3198 = ~( N3127 | N3064 );
	assign N3243 = ~( N3124 | N3193 );
	assign N3404 = ~( N3353 | N3350 );
	assign N3466 = ~( N3404 | N3350 );
	assign N3531 = ~( N3401 | N3461 );
	assign N3693 = ~( N3650 | N3647 );
	assign N3747 = ~( N3693 | N3647 );
	assign N3804 = ~( N3690 | N3742 );
	assign N3992 = ~( N3935 | N3932 );
	assign N4039 = ~( N3992 | N3932 );
	assign N4089 = ~( N3989 | N4034 );
	assign N4281 = ~( N4229 | N4226 );
	assign N4340 = ~( N4281 | N4226 );
	assign N4384 = ~( N4278 | N4335 );
	assign N4578 = ~( N4512 | N4509 );
	assign N4633 = ~( N4578 | N4509 );
	assign N4687 = ~( N4575 | N4628 );
	assign N4866 = ~( N4805 | N4802 );
	assign N4933 = ~( N4866 | N4802 );
	assign N4984 = ~( N4863 | N4928 );
	assign N5163 = ~( N5106 | N5103 );
	assign N5226 = ~( N5163 | N5103 );
	assign N5287 = ~( N5160 | N5221 );
	assign N5467 = ~( N5413 | N5410 );
	assign N5527 = ~( N5467 | N5410 );
	assign N5585 = ~( N5464 | N5522 );
	assign N5776 = ~( N5718 | N5715 );
	assign N5830 = ~( N5776 | N5715 );
	assign N5877 = ~( N5773 | N5825 );
	assign N1676 = ~( N1618 | N1566 );
	assign N1711 = ~( N1676 | N1566 );
	assign N1708 = ~( N1615 | N1672 );
	assign N1995 = ~( N1938 | N1886 );
	assign N2029 = ~( N1995 | N1886 );
	assign N2026 = ~( N1935 | N1991 );
	assign N2260 = ~( N2214 | N2211 );
	assign N2318 = ~( N2260 | N2211 );
	assign N2348 = ~( N2257 | N2313 );
	assign N2539 = ~( N2467 | N2464 );
	assign N2587 = ~( N2539 | N2464 );
	assign N2639 = ~( N2536 | N2582 );
	assign N2797 = ~( N2736 | N2733 );
	assign N2869 = ~( N2797 | N2733 );
	assign N2912 = ~( N2794 | N2864 );
	assign N3070 = ~( N3019 | N3016 );
	assign N3132 = ~( N3070 | N3016 );
	assign N3197 = ~( N3067 | N3127 );
	assign N3356 = ~( N3314 | N3311 );
	assign N3409 = ~( N3356 | N3311 );
	assign N3465 = ~( N3353 | N3404 );
	assign N3653 = ~( N3595 | N3592 );
	assign N3698 = ~( N3653 | N3592 );
	assign N3746 = ~( N3650 | N3693 );
	assign N3938 = ~( N3886 | N3883 );
	assign N3997 = ~( N3938 | N3883 );
	assign N4038 = ~( N3935 | N3992 );
	assign N4232 = ~( N4164 | N4161 );
	assign N4286 = ~( N4232 | N4161 );
	assign N4339 = ~( N4229 | N4281 );
	assign N4515 = ~( N4453 | N4450 );
	assign N4583 = ~( N4515 | N4450 );
	assign N4632 = ~( N4512 | N4578 );
	assign N4808 = ~( N4751 | N4748 );
	assign N4871 = ~( N4808 | N4748 );
	assign N4932 = ~( N4805 | N4866 );
	assign N5109 = ~( N5056 | N5053 );
	assign N5168 = ~( N5109 | N5053 );
	assign N5225 = ~( N5106 | N5163 );
	assign N5416 = ~( N5357 | N5354 );
	assign N5472 = ~( N5416 | N5354 );
	assign N5526 = ~( N5413 | N5467 );
	assign N5721 = ~( N5663 | N5660 );
	assign N5781 = ~( N5721 | N5660 );
	assign N5829 = ~( N5718 | N5776 );
	assign N1680 = ~( N1621 | N1571 );
	assign N1713 = ~( N1680 | N1571 );
	assign N1710 = ~( N1618 | N1676 );
	assign N1941 = ~( N1894 | N1891 );
	assign N2000 = ~( N1941 | N1891 );
	assign N2028 = ~( N1938 | N1995 );
	assign N2217 = ~( N2142 | N2139 );
	assign N2265 = ~( N2217 | N2139 );
	assign N2317 = ~( N2214 | N2260 );
	assign N2470 = ~( N2407 | N2404 );
	assign N2544 = ~( N2470 | N2404 );
	assign N2586 = ~( N2467 | N2539 );
	assign N2739 = ~( N2687 | N2684 );
	assign N2802 = ~( N2739 | N2684 );
	assign N2868 = ~( N2736 | N2797 );
	assign N3022 = ~( N2980 | N2977 );
	assign N3075 = ~( N3022 | N2977 );
	assign N3131 = ~( N3019 | N3070 );
	assign N3317 = ~( N3257 | N3254 );
	assign N3361 = ~( N3317 | N3254 );
	assign N3408 = ~( N3314 | N3356 );
	assign N3598 = ~( N3545 | N3542 );
	assign N3658 = ~( N3598 | N3542 );
	assign N3697 = ~( N3595 | N3653 );
	assign N3889 = ~( N3818 | N3815 );
	assign N3943 = ~( N3889 | N3815 );
	assign N3996 = ~( N3886 | N3938 );
	assign N4167 = ~( N4103 | N4100 );
	assign N4237 = ~( N4167 | N4100 );
	assign N4285 = ~( N4164 | N4232 );
	assign N4456 = ~( N4398 | N4395 );
	assign N4520 = ~( N4456 | N4395 );
	assign N4582 = ~( N4453 | N4515 );
	assign N4754 = ~( N4701 | N4698 );
	assign N4813 = ~( N4754 | N4698 );
	assign N4870 = ~( N4751 | N4808 );
	assign N5059 = ~( N4998 | N4995 );
	assign N5114 = ~( N5059 | N4995 );
	assign N5167 = ~( N5056 | N5109 );
	assign N5360 = ~( N5301 | N5298 );
	assign N5421 = ~( N5360 | N5298 );
	assign N5471 = ~( N5357 | N5416 );
	assign N5666 = ~( N5599 | N5596 );
	assign N5726 = ~( N5666 | N5596 );
	assign N5780 = ~( N5663 | N5721 );
	assign N1712 = ~( N1621 | N1680 );
	assign N1999 = ~( N1894 | N1941 );
	assign N2264 = ~( N2142 | N2217 );
	assign N2543 = ~( N2407 | N2470 );
	assign N2801 = ~( N2687 | N2739 );
	assign N3074 = ~( N2980 | N3022 );
	assign N3360 = ~( N3257 | N3317 );
	assign N3657 = ~( N3545 | N3598 );
	assign N3942 = ~( N3818 | N3889 );
	assign N4236 = ~( N4103 | N4167 );
	assign N4519 = ~( N4398 | N4456 );
	assign N4812 = ~( N4701 | N4754 );
	assign N5113 = ~( N4998 | N5059 );
	assign N5420 = ~( N5301 | N5360 );
	assign N5725 = ~( N5599 | N5666 );
	assign N6281 = ~( N5727 | N6277 );
	assign N6285 = ~( N5727 | N6281 );
	assign N1717 = ~( N1686 | N1687 );
	assign N2037 = ~( N2004 | N2005 );
	assign N2362 = ~( N2326 | N2327 );
	assign N2694 = ~( N2653 | N2654 );
	assign N3028 = ~( N2987 | N2988 );
	assign N3365 = ~( N3323 | N3324 );
	assign N3706 = ~( N3662 | N3663 );
	assign N4052 = ~( N4005 | N4006 );
	assign N4405 = ~( N4353 | N4354 );
	assign N4760 = ~( N4708 | N4709 );
	assign N5118 = ~( N5065 | N5066 );
	assign N5480 = ~( N5425 | N5426 );
	assign N5834 = ~( N5785 | N5786 );
	assign N6061 = ~( N6035 | N6036 );
	assign N6147 = ~( N6124 | N6150 );
	assign N6138 = ~( N6133 | N6134 );
	assign N1720 = ~( N1688 | N1689 );
	assign N2040 = ~( N2006 | N2007 );
	assign N2365 = ~( N2328 | N2329 );
	assign N2697 = ~( N2655 | N2656 );
	assign N3031 = ~( N2989 | N2990 );
	assign N3368 = ~( N3325 | N3326 );
	assign N3709 = ~( N3664 | N3665 );
	assign N4055 = ~( N4007 | N4008 );
	assign N4408 = ~( N4355 | N4356 );
	assign N4763 = ~( N4710 | N4711 );
	assign N5121 = ~( N5067 | N5068 );
	assign N5483 = ~( N5427 | N5428 );
	assign N5837 = ~( N5787 | N5788 );
	assign N6037 = ~( N6009 | N6010 );
	assign N6157 = ~( N6114 | N6151 );
	assign N6135 = ~( N6128 | N6129 );
	assign N1723 = ~( N1690 | N1691 );
	assign N2043 = ~( N2008 | N2009 );
	assign N2368 = ~( N2330 | N2331 );
	assign N2700 = ~( N2657 | N2658 );
	assign N3034 = ~( N2991 | N2992 );
	assign N3371 = ~( N3327 | N3328 );
	assign N3712 = ~( N3666 | N3667 );
	assign N4058 = ~( N4009 | N4010 );
	assign N4411 = ~( N4357 | N4358 );
	assign N4766 = ~( N4712 | N4713 );
	assign N5124 = ~( N5069 | N5070 );
	assign N5486 = ~( N5429 | N5430 );
	assign N5789 = ~( N5738 | N5739 );
	assign N6011 = ~( N5979 | N5980 );
	assign N6167 = ~( N6097 | N6161 );
	assign N6130 = ~( N6118 | N6119 );
	assign N1726 = ~( N1692 | N1693 );
	assign N2046 = ~( N2010 | N2011 );
	assign N2371 = ~( N2332 | N2333 );
	assign N2703 = ~( N2659 | N2660 );
	assign N3037 = ~( N2993 | N2994 );
	assign N3374 = ~( N3329 | N3330 );
	assign N3715 = ~( N3668 | N3669 );
	assign N4061 = ~( N4011 | N4012 );
	assign N4414 = ~( N4359 | N4360 );
	assign N4769 = ~( N4714 | N4715 );
	assign N5127 = ~( N5071 | N5072 );
	assign N5431 = ~( N5378 | N5379 );
	assign N5740 = ~( N5683 | N5684 );
	assign N5981 = ~( N5945 | N5946 );
	assign N6177 = ~( N6076 | N6171 );
	assign N6120 = ~( N6101 | N6102 );
	assign N1729 = ~( N1694 | N1695 );
	assign N2049 = ~( N2012 | N2013 );
	assign N2374 = ~( N2334 | N2335 );
	assign N2706 = ~( N2661 | N2662 );
	assign N3040 = ~( N2995 | N2996 );
	assign N3377 = ~( N3331 | N3332 );
	assign N3718 = ~( N3670 | N3671 );
	assign N4064 = ~( N4013 | N4014 );
	assign N4417 = ~( N4361 | N4362 );
	assign N4772 = ~( N4716 | N4717 );
	assign N5073 = ~( N5021 | N5022 );
	assign N5380 = ~( N5322 | N5323 );
	assign N5685 = ~( N5628 | N5629 );
	assign N5947 = ~( N5902 | N5903 );
	assign N6187 = ~( N6052 | N6181 );
	assign N6103 = ~( N6080 | N6081 );
	assign N1732 = ~( N1696 | N1697 );
	assign N2052 = ~( N2014 | N2015 );
	assign N2377 = ~( N2336 | N2337 );
	assign N2709 = ~( N2663 | N2664 );
	assign N3043 = ~( N2997 | N2998 );
	assign N3380 = ~( N3333 | N3334 );
	assign N3721 = ~( N3672 | N3673 );
	assign N4067 = ~( N4015 | N4016 );
	assign N4420 = ~( N4363 | N4364 );
	assign N4718 = ~( N4666 | N4667 );
	assign N5023 = ~( N4963 | N4964 );
	assign N5324 = ~( N5266 | N5267 );
	assign N5630 = ~( N5564 | N5565 );
	assign N5904 = ~( N5856 | N5857 );
	assign N6197 = ~( N6026 | N6191 );
	assign N6082 = ~( N6056 | N6057 );
	assign N1735 = ~( N1698 | N1699 );
	assign N2055 = ~( N2016 | N2017 );
	assign N2380 = ~( N2338 | N2339 );
	assign N2712 = ~( N2665 | N2666 );
	assign N3046 = ~( N2999 | N3000 );
	assign N3383 = ~( N3335 | N3336 );
	assign N3724 = ~( N3674 | N3675 );
	assign N4070 = ~( N4017 | N4018 );
	assign N4365 = ~( N4318 | N4319 );
	assign N4668 = ~( N4611 | N4612 );
	assign N4965 = ~( N4911 | N4912 );
	assign N5268 = ~( N5204 | N5205 );
	assign N5566 = ~( N5505 | N5506 );
	assign N5858 = ~( N5808 | N5809 );
	assign N6207 = ~( N5996 | N6201 );
	assign N6058 = ~( N6030 | N6031 );
	assign N1738 = ~( N1700 | N1701 );
	assign N2058 = ~( N2018 | N2019 );
	assign N2383 = ~( N2340 | N2341 );
	assign N2715 = ~( N2667 | N2668 );
	assign N3049 = ~( N3001 | N3002 );
	assign N3386 = ~( N3337 | N3338 );
	assign N3727 = ~( N3676 | N3677 );
	assign N4019 = ~( N3975 | N3976 );
	assign N4320 = ~( N4264 | N4265 );
	assign N4613 = ~( N4561 | N4562 );
	assign N4913 = ~( N4849 | N4850 );
	assign N5206 = ~( N5146 | N5147 );
	assign N5507 = ~( N5450 | N5451 );
	assign N5810 = ~( N5759 | N5760 );
	assign N6217 = ~( N5962 | N6211 );
	assign N6032 = ~( N6000 | N6001 );
	assign N1741 = ~( N1702 | N1703 );
	assign N2061 = ~( N2020 | N2021 );
	assign N2386 = ~( N2342 | N2343 );
	assign N2718 = ~( N2669 | N2670 );
	assign N3052 = ~( N3003 | N3004 );
	assign N3389 = ~( N3339 | N3340 );
	assign N3678 = ~( N3636 | N3637 );
	assign N3977 = ~( N3921 | N3922 );
	assign N4266 = ~( N4215 | N4216 );
	assign N4563 = ~( N4498 | N4499 );
	assign N4851 = ~( N4791 | N4792 );
	assign N5148 = ~( N5092 | N5093 );
	assign N5452 = ~( N5399 | N5400 );
	assign N5761 = ~( N5704 | N5705 );
	assign N6227 = ~( N5919 | N6221 );
	assign N6002 = ~( N5966 | N5967 );
	assign N1744 = ~( N1704 | N1705 );
	assign N2064 = ~( N2022 | N2023 );
	assign N2389 = ~( N2344 | N2345 );
	assign N2721 = ~( N2671 | N2672 );
	assign N3055 = ~( N3005 | N3006 );
	assign N3341 = ~( N3300 | N3301 );
	assign N3638 = ~( N3581 | N3582 );
	assign N3923 = ~( N3872 | N3873 );
	assign N4217 = ~( N4150 | N4151 );
	assign N4500 = ~( N4439 | N4440 );
	assign N4793 = ~( N4737 | N4738 );
	assign N5094 = ~( N5042 | N5043 );
	assign N5401 = ~( N5343 | N5344 );
	assign N5706 = ~( N5649 | N5650 );
	assign N6237 = ~( N5873 | N6231 );
	assign N5968 = ~( N5923 | N5924 );
	assign N1747 = ~( N1706 | N1707 );
	assign N2067 = ~( N2024 | N2025 );
	assign N2392 = ~( N2346 | N2347 );
	assign N2724 = ~( N2673 | N2674 );
	assign N3007 = ~( N2966 | N2967 );
	assign N3302 = ~( N3243 | N3244 );
	assign N3583 = ~( N3531 | N3532 );
	assign N3874 = ~( N3804 | N3805 );
	assign N4152 = ~( N4089 | N4090 );
	assign N4441 = ~( N4384 | N4385 );
	assign N4739 = ~( N4687 | N4688 );
	assign N5044 = ~( N4984 | N4985 );
	assign N5345 = ~( N5287 | N5288 );
	assign N5651 = ~( N5585 | N5586 );
	assign N6247 = ~( N5825 | N6241 );
	assign N5925 = ~( N5877 | N5878 );
	assign N1750 = ~( N1708 | N1709 );
	assign N2070 = ~( N2026 | N2027 );
	assign N2395 = ~( N2348 | N2349 );
	assign N2675 = ~( N2639 | N2640 );
	assign N2968 = ~( N2912 | N2913 );
	assign N3245 = ~( N3197 | N3198 );
	assign N3533 = ~( N3465 | N3466 );
	assign N3806 = ~( N3746 | N3747 );
	assign N4091 = ~( N4038 | N4039 );
	assign N4386 = ~( N4339 | N4340 );
	assign N4689 = ~( N4632 | N4633 );
	assign N4986 = ~( N4932 | N4933 );
	assign N5289 = ~( N5225 | N5226 );
	assign N5587 = ~( N5526 | N5527 );
	assign N6257 = ~( N5776 | N6251 );
	assign N5879 = ~( N5829 | N5830 );
	assign N1753 = ~( N1710 | N1711 );
	assign N2073 = ~( N2028 | N2029 );
	assign N2350 = ~( N2317 | N2318 );
	assign N2641 = ~( N2586 | N2587 );
	assign N2914 = ~( N2868 | N2869 );
	assign N3199 = ~( N3131 | N3132 );
	assign N3467 = ~( N3408 | N3409 );
	assign N3748 = ~( N3697 | N3698 );
	assign N4040 = ~( N3996 | N3997 );
	assign N4341 = ~( N4285 | N4286 );
	assign N4634 = ~( N4582 | N4583 );
	assign N4934 = ~( N4870 | N4871 );
	assign N5227 = ~( N5167 | N5168 );
	assign N5528 = ~( N5471 | N5472 );
	assign N6267 = ~( N5721 | N6261 );
	assign N5831 = ~( N5780 | N5781 );
	assign N1756 = ~( N1712 | N1713 );
	assign N2030 = ~( N1999 | N2000 );
	assign N2319 = ~( N2264 | N2265 );
	assign N2588 = ~( N2543 | N2544 );
	assign N2870 = ~( N2801 | N2802 );
	assign N3133 = ~( N3074 | N3075 );
	assign N3410 = ~( N3360 | N3361 );
	assign N3699 = ~( N3657 | N3658 );
	assign N3998 = ~( N3942 | N3943 );
	assign N4287 = ~( N4236 | N4237 );
	assign N4584 = ~( N4519 | N4520 );
	assign N4872 = ~( N4812 | N4813 );
	assign N5169 = ~( N5113 | N5114 );
	assign N5473 = ~( N5420 | N5421 );
	assign N6277 = ~( N5666 | N6271 );
	assign N5782 = ~( N5725 | N5726 );
	assign N6286 = ~( N6281 | N6277 );
	assign N6288 = ~( N6285 | N6286 );
	assign N6151 = ~( N6135 | N6147 );
	assign N6156 = ~( N6151 | N6147 );
	assign N6150 = ~N6138;
	assign N6161 = ~( N6130 | N6157 );
	assign N6166 = ~( N6161 | N6157 );
	assign N6155 = ~( N6135 | N6151 );
	assign N6171 = ~( N6120 | N6167 );
	assign N6176 = ~( N6171 | N6167 );
	assign N6165 = ~( N6130 | N6161 );
	assign N6181 = ~( N6103 | N6177 );
	assign N6186 = ~( N6181 | N6177 );
	assign N6175 = ~( N6120 | N6171 );
	assign N6191 = ~( N6082 | N6187 );
	assign N6196 = ~( N6191 | N6187 );
	assign N6185 = ~( N6103 | N6181 );
	assign N6201 = ~( N6058 | N6197 );
	assign N6206 = ~( N6201 | N6197 );
	assign N6195 = ~( N6082 | N6191 );
	assign N6211 = ~( N6032 | N6207 );
	assign N6216 = ~( N6211 | N6207 );
	assign N6205 = ~( N6058 | N6201 );
	assign N6221 = ~( N6002 | N6217 );
	assign N6226 = ~( N6221 | N6217 );
	assign N6215 = ~( N6032 | N6211 );
	assign N6231 = ~( N5968 | N6227 );
	assign N6236 = ~( N6231 | N6227 );
	assign N6225 = ~( N6002 | N6221 );
	assign N6241 = ~( N5925 | N6237 );
	assign N6246 = ~( N6241 | N6237 );
	assign N6235 = ~( N5968 | N6231 );
	assign N6251 = ~( N5879 | N6247 );
	assign N6256 = ~( N6251 | N6247 );
	assign N6245 = ~( N5925 | N6241 );
	assign N6261 = ~( N5831 | N6257 );
	assign N6266 = ~( N6261 | N6257 );
	assign N6255 = ~( N5879 | N6251 );
	assign N6271 = ~( N5782 | N6267 );
	assign N6276 = ~( N6271 | N6267 );
	assign N6265 = ~( N5831 | N6261 );
	assign N6275 = ~( N5782 | N6271 );
	assign N6160 = ~( N6155 | N6156 );
	assign N6170 = ~( N6165 | N6166 );
	assign N6180 = ~( N6175 | N6176 );
	assign N6190 = ~( N6185 | N6186 );
	assign N6200 = ~( N6195 | N6196 );
	assign N6210 = ~( N6205 | N6206 );
	assign N6220 = ~( N6215 | N6216 );
	assign N6230 = ~( N6225 | N6226 );
	assign N6240 = ~( N6235 | N6236 );
	assign N6250 = ~( N6245 | N6246 );
	assign N6260 = ~( N6255 | N6256 );
	assign N6270 = ~( N6265 | N6266 );
	assign N6280 = ~( N6275 | N6276 );
endmodule
