module c499(N135, N133, N136, N132, N129, N121, N117, N9, N37, N45, N77, N33, N29, N25, N49, N134, N13, N131, N41, N21, N57, N5, N61, N17, N69, N137, N85, N1, N125, N53, N73, N101, N130, N113, N65, N81, N89, N109, N105, N93, N97, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, N755, N753, N725, N734, N750, N754, N736, N741, N747, N730, N735, N728, N744, N748, N732, N727, N726, N724, N737, N731, N738, N733, N739, N749, N729, N740, N742, N751, N743, N745, N746, N752);
	input N135, N133, N136, N132, N129, N121, N117, N9, N37, N45, N77, N33, N29, N25, N49, N134, N13, N131, N41, N21, N57, N5, N61, N17, N69, N137, N85, N1, N125, N53, N73, N101, N130, N113, N65, N81, N89, N109, N105, N93, N97;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9;
	output N755, N753, N725, N734, N750, N754, N736, N741, N747, N730, N735, N728, N744, N748, N732, N727, N726, N724, N737, N731, N738, N733, N739, N749, N729, N740, N742, N751, N743, N745, N746, N752;
	wire N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N250, N274, N724, N276, N725, N251, N278, N726, N280, N727, N252, N728, N729, N253, N730, N731, N254, N275, N732, N277, N733, N255, N279, N734, N281, N735, N256, N736, N737, N257, N738, N739, N258, N282, N740, N284, N741, N259, N286, N742, N288, N743, N260, N744, N745, N261, N746, N747, N262, N283, N748, N285, N749, N263, N287, N750, N289, N751, N264, N752, N753, N265, N754, N755, N266, N267, N268, N269, N270, N271, N272, N273, N290, N314, N315, N316, N317, N293, N296, N299, N302, N318, N319, N320, N321, N305, N308, N311, N346, N347, N348, N349, N350, N351, N352, N353, N338, N340, N354, N367, N380, N393, N341, N339, N342, N344, N406, N419, N432, N445, N345, N343, N692, N696, N700, N704, N597, N554, n_78, N693, N697, N701, N705, N596, N555, n_80, N694, N698, N702, N706, N595, N556, N640, N650, N695, N699, N703, N707, N594, N559, N645, N655, N708, N712, N716, N720, N601, N570, n_74, N709, N713, N717, N721, N600, N566, n_76, N710, N714, N718, N722, N599, N569, N620, N630, N711, N715, N719, N723, N598, N567, N625, N635, N602, N607;
	wire N607_key, N602_key, N597_key, N596_key, N595_key, N594_key, N601_key, N600_key, N599_key, N598_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9;
	assign N250 = ( N1 ^ N5 );
	assign N274 = ( N1 ^ N17 );
	assign N724 = ( N1 ^ N692 );
	assign N276 = ( N5 ^ N21 );
	assign N725 = ( N5 ^ N693 );
	assign N251 = ( N9 ^ N13 );
	assign N278 = ( N9 ^ N25 );
	assign N726 = ( N9 ^ N694 );
	assign N280 = ( N13 ^ N29 );
	assign N727 = ( N13 ^ N695 );
	assign N252 = ( N17 ^ N21 );
	assign N728 = ( N17 ^ N696 );
	assign N729 = ( N21 ^ N697 );
	assign N253 = ( N25 ^ N29 );
	assign N730 = ( N25 ^ N698 );
	assign N731 = ( N29 ^ N699 );
	assign N254 = ( N33 ^ N37 );
	assign N275 = ( N33 ^ N49 );
	assign N732 = ( N33 ^ N700 );
	assign N277 = ( N37 ^ N53 );
	assign N733 = ( N37 ^ N701 );
	assign N255 = ( N41 ^ N45 );
	assign N279 = ( N41 ^ N57 );
	assign N734 = ( N41 ^ N702 );
	assign N281 = ( N45 ^ N61 );
	assign N735 = ( N45 ^ N703 );
	assign N256 = ( N49 ^ N53 );
	assign N736 = ( N49 ^ N704 );
	assign N737 = ( N53 ^ N705 );
	assign N257 = ( N57 ^ N61 );
	assign N738 = ( N57 ^ N706 );
	assign N739 = ( N61 ^ N707 );
	assign N258 = ( N65 ^ N69 );
	assign N282 = ( N65 ^ N81 );
	assign N740 = ( N65 ^ N708 );
	assign N284 = ( N69 ^ N85 );
	assign N741 = ( N69 ^ N709 );
	assign N259 = ( N73 ^ N77 );
	assign N286 = ( N73 ^ N89 );
	assign N742 = ( N73 ^ N710 );
	assign N288 = ( N77 ^ N93 );
	assign N743 = ( N77 ^ N711 );
	assign N260 = ( N81 ^ N85 );
	assign N744 = ( N81 ^ N712 );
	assign N745 = ( N85 ^ N713 );
	assign N261 = ( N89 ^ N93 );
	assign N746 = ( N89 ^ N714 );
	assign N747 = ( N93 ^ N715 );
	assign N262 = ( N97 ^ N101 );
	assign N283 = ( N97 ^ N113 );
	assign N748 = ( N97 ^ N716 );
	assign N285 = ( N101 ^ N117 );
	assign N749 = ( N101 ^ N717 );
	assign N263 = ( N105 ^ N109 );
	assign N287 = ( N105 ^ N121 );
	assign N750 = ( N105 ^ N718 );
	assign N289 = ( N109 ^ N125 );
	assign N751 = ( N109 ^ N719 );
	assign N264 = ( N113 ^ N117 );
	assign N752 = ( N113 ^ N720 );
	assign N753 = ( N117 ^ N721 );
	assign N265 = ( N121 ^ N125 );
	assign N754 = ( N121 ^ N722 );
	assign N755 = ( N125 ^ N723 );
	assign N266 = ( N129 & N137 );
	assign N267 = ( N130 & N137 );
	assign N268 = ( N131 & N137 );
	assign N269 = ( N132 & N137 );
	assign N270 = ( N133 & N137 );
	assign N271 = ( N134 & N137 );
	assign N272 = ( N135 & N137 );
	assign N273 = ( N136 & N137 );
	assign N290 = ( N250 ^ N251 );
	assign N314 = ( N274 ^ N275 );
	assign N315 = ( N276 ^ N277 );
	assign N316 = ( N278 ^ N279 );
	assign N317 = ( N280 ^ N281 );
	assign N293 = ( N252 ^ N253 );
	assign N296 = ( N254 ^ N255 );
	assign N299 = ( N256 ^ N257 );
	assign N302 = ( N258 ^ N259 );
	assign N318 = ( N282 ^ N283 );
	assign N319 = ( N284 ^ N285 );
	assign N320 = ( N286 ^ N287 );
	assign N321 = ( N288 ^ N289 );
	assign N305 = ( N260 ^ N261 );
	assign N308 = ( N262 ^ N263 );
	assign N311 = ( N264 ^ N265 );
	assign N346 = ( N266 ^ N342 );
	assign N347 = ( N267 ^ N343 );
	assign N348 = ( N268 ^ N344 );
	assign N349 = ( N269 ^ N345 );
	assign N350 = ( N270 ^ N338 );
	assign N351 = ( N271 ^ N339 );
	assign N352 = ( N272 ^ N340 );
	assign N353 = ( N273 ^ N341 );
	assign N338 = ( N290 ^ N293 );
	assign N340 = ( N290 ^ N296 );
	assign N354 = ( N314 ^ N346 );
	assign N367 = ( N315 ^ N347 );
	assign N380 = ( N316 ^ N348 );
	assign N393 = ( N317 ^ N349 );
	assign N341 = ( N293 ^ N299 );
	assign N339 = ( N296 ^ N299 );
	assign N342 = ( N302 ^ N305 );
	assign N344 = ( N302 ^ N308 );
	assign N406 = ( N318 ^ N350 );
	assign N419 = ( N319 ^ N351 );
	assign N432 = ( N320 ^ N352 );
	assign N445 = ( N321 ^ N353 );
	assign N345 = ( N305 ^ N311 );
	assign N343 = ( N308 ^ N311 );
	assign N692 = ( N354 & N620 );
	assign N696 = ( N354 & N625 );
	assign N700 = ( N354 & N630 );
	assign N704 = ( N354 & N635 );
	assign N597 = ( N354 & N555 & N556 & N559 );
	assign N554 = ~N354;
	assign n_78 = ( N354 & N555 );
	assign N693 = ( N367 & N620 );
	assign N697 = ( N367 & N625 );
	assign N701 = ( N367 & N630 );
	assign N705 = ( N367 & N635 );
	assign N596 = ( N554 & N367 & N556 & N559 );
	assign N555 = ~N367;
	assign n_80 = ( N554 & N367 );
	assign N694 = ( N380 & N620 );
	assign N698 = ( N380 & N625 );
	assign N702 = ( N380 & N630 );
	assign N706 = ( N380 & N635 );
	assign N595 = ( N554 & N555 & N380 & N559 );
	assign N556 = ~N380;
	assign N640 = ( N380 & N559 & N607_key & n_78 );
	assign N650 = ( N380 & N559 & N607_key & n_80 );
	assign N695 = ( N393 & N620 );
	assign N699 = ( N393 & N625 );
	assign N703 = ( N393 & N630 );
	assign N707 = ( N393 & N635 );
	assign N594 = ( N554 & N555 & N556 & N393 );
	assign N559 = ~N393;
	assign N645 = ( N556 & N393 & N607_key & n_78 );
	assign N655 = ( N556 & N393 & N607_key & n_80 );
	assign N708 = ( N406 & N640 );
	assign N712 = ( N406 & N645 );
	assign N716 = ( N406 & N650 );
	assign N720 = ( N406 & N655 );
	assign N601 = ( N406 & N566 & N569 & N567 );
	assign N570 = ~N406;
	assign n_74 = ( N406 & N566 );
	assign N709 = ( N419 & N640 );
	assign N713 = ( N419 & N645 );
	assign N717 = ( N419 & N650 );
	assign N721 = ( N419 & N655 );
	assign N600 = ( N570 & N419 & N569 & N567 );
	assign N566 = ~N419;
	assign n_76 = ( N570 & N419 );
	assign N710 = ( N432 & N640 );
	assign N714 = ( N432 & N645 );
	assign N718 = ( N432 & N650 );
	assign N722 = ( N432 & N655 );
	assign N599 = ( N570 & N566 & N432 & N567 );
	assign N569 = ~N432;
	assign N620 = ( N432 & N567 & N602_key & n_74 );
	assign N630 = ( N432 & N567 & N602_key & n_76 );
	assign N711 = ( N445 & N640 );
	assign N715 = ( N445 & N645 );
	assign N719 = ( N445 & N650 );
	assign N723 = ( N445 & N655 );
	assign N598 = ( N570 & N566 & N569 & N445 );
	assign N567 = ~N445;
	assign N625 = ( N569 & N445 & N602_key & n_74 );
	assign N635 = ( N569 & N445 & N602_key & n_76 );
	assign N602 = ( N594_key | N595_key | N596_key | N597_key );
	assign N607 = ( N598_key | N599_key | N600_key | N601_key );
	assign N607_key = ~( N607 ^ key_0 );
	assign N602_key = ~( N602 ^ key_1 );
	assign N597_key = ~( N597 ^ key_2 );
	assign N596_key = ~( N596 ^ key_3 );
	assign N595_key = ~( N595 ^ key_4 );
	assign N594_key = ~( N594 ^ key_5 );
	assign N601_key = ~( N601 ^ key_6 );
	assign N600_key = ~( N600 ^ key_7 );
	assign N599_key = ~( N599 ^ key_8 );
	assign N598_key = ~( N598 ^ key_9 );
endmodule
