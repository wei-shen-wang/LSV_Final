module c432(N115, N112, N108, N102, N27, N24, N21, N11, N37, N30, N95, N56, N8, N99, N1, N92, N63, N4, N43, N40, N50, N34, N53, N60, N82, N17, N69, N14, N47, N73, N105, N86, N76, N79, N66, N89, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, N431, N430, N432, N421, N370, N329, N223);
	input N115, N112, N108, N102, N27, N24, N21, N11, N37, N30, N95, N56, N8, N99, N1, N92, N63, N4, N43, N40, N50, N34, N53, N60, N82, N17, N69, N14, N47, N73, N105, N86, N76, N79, N66, N89;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9;
	output N431, N430, N432, N421, N370, N329, N223;
	wire N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N242, N118, N154, N380, N119, N334, N157, N246, N122, N371, N158, N159, N381, N123, N336, N183, N250, N126, N372, N184, N162, N386, N127, N338, N185, N254, N130, N373, N186, N165, N393, N131, N340, N187, N255, N134, N374, N188, N168, N399, N135, N342, N189, N256, N138, N375, N190, N171, N404, N139, N344, N191, N257, N142, N376, N192, N174, N407, N143, N345, N193, N258, N146, N377, N194, N177, N411, N147, N346, N195, N259, N150, N378, N196, N180, N414, N151, N347, N197, N379, N198, N224, n_44, N415, N260, N263, N227, N430, N431, N432, n_56, N264, N288, N230, N422, N425, N429, N267, N289, N233, n_45, N428, N417, n_57, N270, N290, N236, N273, N291, N239, n_46, N418, n_58, N276, N292, N243, N419, N279, N293, N247, n_47, N420, n_59, N282, N294, N251, N285, N295, N199, N421, N330, n_48, N300, N416, N331, N301, N332, N302, N333, n_49, N303, N335, N304, N337, n_50, N305, N339, N306, N341, n_51, N307, N343, N308, N223, N348, N296, N349, N350, N351, N352, N353, N354, N355, N356, n_52, N329, n_53, n_54, n_55, N357, N370;
	wire N357_key, n_55_key, N14_key, N27_key, N40_key, N53_key, N66_key, N79_key, N92_key, N105_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9;
	assign N242 = ~( N1 & N223 );
	assign N118 = ~N1;
	assign N154 = ~( N118 & N4 );
	assign N380 = ~( N4 & N242 & N334 & N371 );
	assign N119 = ~N4;
	assign N334 = ~( N8 & N329 );
	assign N157 = ~( N8 | N119 );
	assign N246 = ~( N223 & N11 );
	assign N122 = ~N11;
	assign N371 = ~( N14_key & N370 );
	assign N158 = ~( N14_key | N119 );
	assign N159 = ~( N122 & N17 );
	assign N381 = ~( N246 & N336 & N372 & N17 );
	assign N123 = ~N17;
	assign N336 = ~( N329 & N21 );
	assign N183 = ~( N21 | N123 );
	assign N250 = ~( N223 & N24 );
	assign N126 = ~N24;
	assign N372 = ~( N370 & N27_key );
	assign N184 = ~( N27_key | N123 );
	assign N162 = ~( N126 & N30 );
	assign N386 = ~( N250 & N338 & N373 & N30 );
	assign N127 = ~N30;
	assign N338 = ~( N329 & N34 );
	assign N185 = ~( N34 | N127 );
	assign N254 = ~( N223 & N37 );
	assign N130 = ~N37;
	assign N373 = ~( N370 & N40_key );
	assign N186 = ~( N40_key | N127 );
	assign N165 = ~( N130 & N43 );
	assign N393 = ~( N254 & N340 & N374 & N43 );
	assign N131 = ~N43;
	assign N340 = ~( N329 & N47 );
	assign N187 = ~( N47 | N131 );
	assign N255 = ~( N223 & N50 );
	assign N134 = ~N50;
	assign N374 = ~( N370 & N53_key );
	assign N188 = ~( N53_key | N131 );
	assign N168 = ~( N134 & N56 );
	assign N399 = ~( N255 & N342 & N375 & N56 );
	assign N135 = ~N56;
	assign N342 = ~( N329 & N60 );
	assign N189 = ~( N60 | N135 );
	assign N256 = ~( N223 & N63 );
	assign N138 = ~N63;
	assign N375 = ~( N370 & N66_key );
	assign N190 = ~( N66_key | N135 );
	assign N171 = ~( N138 & N69 );
	assign N404 = ~( N256 & N344 & N376 & N69 );
	assign N139 = ~N69;
	assign N344 = ~( N329 & N73 );
	assign N191 = ~( N73 | N139 );
	assign N257 = ~( N223 & N76 );
	assign N142 = ~N76;
	assign N376 = ~( N370 & N79_key );
	assign N192 = ~( N79_key | N139 );
	assign N174 = ~( N142 & N82 );
	assign N407 = ~( N257 & N345 & N377 & N82 );
	assign N143 = ~N82;
	assign N345 = ~( N329 & N86 );
	assign N193 = ~( N86 | N143 );
	assign N258 = ~( N223 & N89 );
	assign N146 = ~N89;
	assign N377 = ~( N370 & N92_key );
	assign N194 = ~( N92_key | N143 );
	assign N177 = ~( N146 & N95 );
	assign N411 = ~( N258 & N346 & N378 & N95 );
	assign N147 = ~N95;
	assign N346 = ~( N329 & N99 );
	assign N195 = ~( N99 | N147 );
	assign N259 = ~( N223 & N102 );
	assign N150 = ~N102;
	assign N378 = ~( N370 & N105_key );
	assign N196 = ~( N105_key | N147 );
	assign N180 = ~( N150 & N108 );
	assign N414 = ~( N259 & N347 & N379 & N108 );
	assign N151 = ~N108;
	assign N347 = ~( N329 & N112 );
	assign N197 = ~( N112 | N151 );
	assign N379 = ~( N370 & N115 );
	assign N198 = ~( N115 | N151 );
	assign N224 = ( N223 ^ N154 );
	assign n_44 = ( N154 & N159 & N162 );
	assign N415 = ~N380;
	assign N260 = ~( N224 & N157 );
	assign N263 = ~( N224 & N158 );
	assign N227 = ( N223 ^ N159 );
	assign N430 = ~( N381 & N386 & N422 & N399 );
	assign N431 = ~( N381 & N386 & N425 & N428 );
	assign N432 = ~( N381 & N422 & N425 & N429 );
	assign n_56 = ( N381 & N386 );
	assign N264 = ~( N227 & N183 );
	assign N288 = ~( N227 & N184 );
	assign N230 = ( N223 ^ N162 );
	assign N422 = ~( N386 & N417 );
	assign N425 = ~( N386 & N393 & N418 & N399 );
	assign N429 = ~( N386 & N393 & N407 & N420 );
	assign N267 = ~( N230 & N185 );
	assign N289 = ~( N230 & N186 );
	assign N233 = ( N223 ^ N165 );
	assign n_45 = ( N165 & N168 );
	assign N428 = ~( N399 & N393 & N419 );
	assign N417 = ~N393;
	assign n_57 = ( N393 & N399 );
	assign N270 = ~( N233 & N187 );
	assign N290 = ~( N233 & N188 );
	assign N236 = ( N223 ^ N168 );
	assign N273 = ~( N236 & N189 );
	assign N291 = ~( N236 & N190 );
	assign N239 = ( N223 ^ N171 );
	assign n_46 = ( N171 & N174 );
	assign N418 = ~N404;
	assign n_58 = ( N404 & N407 );
	assign N276 = ~( N239 & N191 );
	assign N292 = ~( N239 & N192 );
	assign N243 = ( N223 ^ N174 );
	assign N419 = ~N407;
	assign N279 = ~( N243 & N193 );
	assign N293 = ~( N243 & N194 );
	assign N247 = ( N223 ^ N177 );
	assign n_47 = ( N177 & N180 );
	assign N420 = ~N411;
	assign n_59 = ( N411 & N414 );
	assign N282 = ~( N247 & N195 );
	assign N294 = ~( N247 & N196 );
	assign N251 = ( N223 ^ N180 );
	assign N285 = ~( N251 & N197 );
	assign N295 = ~( N251 & N198 );
	assign N199 = ( n_44 & n_45 & n_46 & n_47 );
	assign N421 = ~( N415 | N416 );
	assign N330 = ( N329 ^ N260 );
	assign n_48 = ( N260 & N264 & N267 );
	assign N300 = ~N263;
	assign N416 = ( n_56 & n_57 & n_58 & n_59 );
	assign N331 = ( N329 ^ N264 );
	assign N301 = ~N288;
	assign N332 = ( N329 ^ N267 );
	assign N302 = ~N289;
	assign N333 = ( N329 ^ N270 );
	assign n_49 = ( N270 & N273 );
	assign N303 = ~N290;
	assign N335 = ( N329 ^ N273 );
	assign N304 = ~N291;
	assign N337 = ( N329 ^ N276 );
	assign n_50 = ( N276 & N279 );
	assign N305 = ~N292;
	assign N339 = ( N329 ^ N279 );
	assign N306 = ~N293;
	assign N341 = ( N329 ^ N282 );
	assign n_51 = ( N282 & N285 );
	assign N307 = ~N294;
	assign N343 = ( N329 ^ N285 );
	assign N308 = ~N295;
	assign N223 = ~N199;
	assign N348 = ~( N330 & N300 );
	assign N296 = ( n_48 & n_49 & n_50 & n_51 );
	assign N349 = ~( N331 & N301 );
	assign N350 = ~( N332 & N302 );
	assign N351 = ~( N333 & N303 );
	assign N352 = ~( N335 & N304 );
	assign N353 = ~( N337 & N305 );
	assign N354 = ~( N339 & N306 );
	assign N355 = ~( N341 & N307 );
	assign N356 = ~( N343 & N308 );
	assign n_52 = ( N348 & N349 & N350 );
	assign N329 = ~N296;
	assign n_53 = ( N351 & N352 );
	assign n_54 = ( N353 & N354 );
	assign n_55 = ( N355 & N356 );
	assign N357 = ( n_52 & n_53 & n_54 & n_55_key );
	assign N370 = ~N357_key;
	assign N357_key = ~( N357 ^ key_0 );
	assign n_55_key = ~( n_55 ^ key_1 );
	assign N14_key = ~( N14 ^ key_2 );
	assign N27_key = ~( N27 ^ key_3 );
	assign N40_key = ~( N40 ^ key_4 );
	assign N53_key = ~( N53 ^ key_5 );
	assign N66_key = ~( N66 ^ key_6 );
	assign N79_key = ~( N79 ^ key_7 );
	assign N92_key = ~( N92 ^ key_8 );
	assign N105_key = ~( N105 ^ key_9 );
endmodule
