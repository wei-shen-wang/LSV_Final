module cavlc(\trailingones[1], \ctable[2], \ctable[1], \ctable[0], \totalcoeffs[4], \trailingones[0], \totalcoeffs[3], \totalcoeffs[2], \totalcoeffs[1], \totalcoeffs[0], key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, \ctoken_len[4], \ctoken_len[3], \ctoken_len[1], \coeff_token[4], \ctoken_len[2], \coeff_token[3], \ctoken_len[0], \coeff_token[2], \coeff_token[5], \coeff_token[1], \coeff_token[0]);
	input \trailingones[1], \ctable[2], \ctable[1], \ctable[0], \totalcoeffs[4], \trailingones[0], \totalcoeffs[3], \totalcoeffs[2], \totalcoeffs[1], \totalcoeffs[0];
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62;
	output \ctoken_len[4], \ctoken_len[3], \ctoken_len[1], \coeff_token[4], \ctoken_len[2], \coeff_token[3], \ctoken_len[0], \coeff_token[2], \coeff_token[5], \coeff_token[1], \coeff_token[0];
	wire \totalcoeffs[0], \totalcoeffs[1], \totalcoeffs[2], \totalcoeffs[3], \totalcoeffs[4], \ctable[0], \ctable[1], \ctable[2], \trailingones[0], \trailingones[1], n_9, n28, n42, n60, n75, n144, n172, n195, n202, n203, n217, n230, n317, n396, n441, n471, n480, n522, n560, n643, n674, n_6, n25, n30, n37, n45, n55, n56, n77, n105, n185, n206, n225, n265, n275, n283, n304, n320, n345, n371, n390, n414, n501, n539, n577, n632, n687, n_22, n62, n78, n84, n95, n103, n158, n211, n243, n261, n272, n307, n321, n325, n353, n366, n372, n377, n399, n436, n443, n446, n472, n497, n506, n535, n578, n593, n641, n645, n697, n711, n_3, n89, n110, n198, n214, n226, n232, n259, n262, n281, n310, n328, n352, n368, n386, n398, n413, n423, n490, n531, n545, n554, n568, n571, n677, n690, n_99, n127, n132, n293, n515, n603, n669, n691, n_4, n79, n94, n130, n134, n149, n162, n173, n192, n231, n260, n274, n301, n311, n363, n367, n381, n439, n448, n491, n561, n582, n610, n_54, n73, n91, n100, n109, n128, n131, n151, n170, n179, n210, n235, n266, n276, n282, n323, n329, n451, n499, n701, n_16, n51, n249, n457, n464, n675, n_39, n81, n102, n150, n154, n186, n201, n215, n263, n290, n299, n314, n324, n331, n356, n445, n458, n520, n564, n586, n624, n646, n23, n24, n_13, n41, n53, n161, n174, n238, n255, n401, n452, n484, n525, n636, n36, n63, n70, n74, n98, n107, n116, n153, n200, n298, n376, n425, n442, n461, n474, n485, n543, n546, n562, n570, n594, n609, n654, n142, n_14, n85, n346, n_30, n583, n61, n596, n_59, n343, n145, n462, n_439, n_134, n_153, n_159, n_158, n337, n622, n670, n_169, n479, n_182, n_253, n418, n_364, n_390, n_394, n_437, n_465, n_537, n_619, n29, n44, n82, n108, n139, n169, n197, n212, n216, n227, n271, n279, n362, n406, n435, n509, n553, n585, n640, n659, n699, n296, n_12, n_17, n96, n247, n487, n_26, n627, n_33, n_45, n_44, n92, n_82, n_145, n_162, n_177, n_212, n_219, n284, n_503, n_244, n_265, n660, n_281, n_299, n_321, n415, n_419, n_462, n_489, n_523, n_620, n34, n35, n40, n90, n140, n146, n177, n180, n199, n278, n312, n335, n359, n378, n384, n408, n465, n482, n505, n529, n542, n579, n621, n680, n694, n220, n614, n64, n187, n_258, n459, n_75, n302, n565, n657, n104, n616, n_562, n_122, n_166, n_194, n422, n_207, n_217, n_245, n_256, n_260, n_285, n_297, n_300, n_306, n_325, n681, n_360, n_365, n_368, n_391, n_408, n550, n507, n_543, n_445, n_481, n587, n_531, n_535, n_583, n_595, n22, n67, n191, n193, n309, n383, n391, n469, n530, n536, n567, n676, n684, n692, n121, n_85, n_155, n_171, n228, n_311, n_181, n236, n_206, n_208, n_614, n_247, n633, n_270, n_284, n_296, n_313, n650, n_327, n523, n_350, n431, n710, n_421, n_440, n_458, n556, n574, n_471, n_474, n_563, n_578, n124, n160, n189, n240, n289, n339, n355, n374, n419, n514, n601, n665, n253, n350, n_124, n_105, n_349, n516, n666, n605, n_618, n_577, n52, n57, n72, n87, n115, n222, n292, n342, n478, n559, n625, n682, n700, n_62, n_78, n_108, n_107, \coeff_token[4], \coeff_token[5], n_121, n_125, n175, n_157, n_152, n392, n_180, n_209, n_613, n_239, n_248, n364, n_336, n_294, n382, n_335, n_362, n_371, n492, n607, n_484, n_507, n69, n126, n164, n178, n209, n258, n319, n385, n409, n438, n493, n533, n541, n549, n590, n639, n644, n663, n683, n_61, n_72, n_79, n_84, n_102, n_104, n_115, n_133, n526, n_137, n_165, n_184, n267, n397, n402, n_220, n_432, n555, n_261, n_263, n647, n454, n_411, n_617, n31, n48, n122, n242, n341, \coeff_token[3], n428, n433, n456, n512, n518, n592, n652, n671, n673, n713, n595, n_200, n_377, n50, n83, n113, n117, n125, n136, n155, n246, n404, n496, n502, n573, n619, n695, n708, n_68, n_114, n181, n_117, n_215, n_205, n634, n_170, n678, n688, n_210, n_231, n_237, n315, n_255, n_259, n_267, n357, n_372, n_370, n_378, n_430, n_468, n_567, n_519, n_534, n_11, n71, n_10, n494, n39, n183, n224, n270, n277, n380, n394, n437, n504, n548, n629, n656, n_29, n_42, n_128, n_202, n_188, n_203, n_330, n_374, n_400, n_435, n_527, n_25, n_193, n430, n167, n_58, n147, n99, n_514, n_88, n118, n_119, n_161, n_276, n_346, n426, n_355, n667, n_383, n476, n_413, n_399, n_451, n_453, n_466, n_473, n_495, n_512, n_545, \coeff_token[0], n_66, n_282, n43, n_485, n_48, n_496, n76, n_279, n_111, n_381, n532, n176, n196, n205, n655, n204, n486, n503, n_274, n_516, n_559, n244, n_396, n234, n318, n_345, n444, n473, n481, n547, n528, n563, n649, \ctoken_len[3], n_18, n_32, n_64, n111, n_242, n268, n_148, n_163, n_167, n598, n_610, n_216, n_223, n_302, n_359, n_420, n_460, n_487, n_530, n_550, n_234, n26, n709, n330, n_76, n_197, n_401, n38, n_520, n46, n256, n59, n58, n_73, n106, n188, n207, n229, n269, n_615, n608, n308, n332, n410, n470, n_551, n347, n373, n395, n510, n558, n589, n635, n_36, n_24, n_28, n_71, n_558, n_542, n_142, n_138, n_156, n_222, n313, n_271, n360, n_307, n_314, n_338, n_384, n_397, n_416, n_447, n_450, n_480, n_515, n_571, n_582, n_172, n_510, n65, n_199, n_146, n453, n569, n_379, n97, n112, n_240, n_469, n_548, n_81, n_511, n159, n213, n245, n_352, n630, n273, n322, n326, n354, n370, n379, n400, n447, n498, n_457, n_417, n653, n537, n581, n_488, n642, n648, n698, n712, n27, n599, n_506, n662, n_52, n_190, n_151, n333, n_252, n_310, n_318, n_423, n_442, n_446, n_478, n_564, n696, n_570, n_579, n_95, n221, n_178, n233, n_185, n631, n288, n336, n369, n387, n_540, n403, n_433, n424, n_357, n511, n552, n_461, n_477, n626, n572, n693, n_130, n_149, n_191, n_233, n_277, n_289, n_303, n_347, n_428, n_501, n_556, \coeff_token[1], \coeff_token[2], n163, n133, n165, n_426, n_502, n_41, n_333, n_57, n_69, n_175, n_612, n467, n_576, \ctoken_len[4], n_402, n_491, n_518, n_569, n_585, n80, n101, n137, n135, n358, n517, n_135, n_319, n264, n303, n_292, n_309, n440, n449, n_405, n_504, n584, n611, n_96, n_101, n_127, n_139, n_174, n_616, n_273, n_312, n411, n_573, n_361, n_404, n_443, n_455, n_492, n_539, n_533, n_554, n_568, n93, n129, n152, n521, n689, n171, n_436, n237, n_295, n_324, n_328, n524, n327, n_536, n_375, n500, n32, n_37, n_97, n_386, n_424, n_429, n_498, n_553, n_560, n_561, n250, n_51, n_65, n_89, n_367, n_236, n_109, n_118, n_196, n_331, n_410, n_414, n_476, n_528, n_581, n_593, n88, n194, n_140, n156, n_524, n_565, n_574, n291, n305, n300, n_250, n334, n_287, n450, n566, n628, n_56, n_406, n_34, n_143, n_187, n_221, n_316, n_322, n_456, n_526, n_547, n54, n166, n540, n239, n257, n405, n488, n527, n637, n_356, n_131, n344, n_112, n620, n114, n157, n340, n420, n_353, n_557, n466, n_392, n544, n597, n618, n86, n_31, n66, n_60, n148, n463, n_441, n_136, n_154, n_160, n_546, n_415, n338, n623, n_195, n483, n_183, n_254, n_366, n477, n_395, n_454, n_438, n_467, n_538, n_86, n306, n_213, n190, n208, n475, n280, n375, n615, n557, n588, n672, n661, n297, n_594, n_264, n460, n248, n_27, n47, n_204, n_47, n_46, n_83, n_147, n_179, n_214, n_505, n_246, n_266, n_337, n_389, n_611, n_301, n_323, n_463, n_490, n_525, n49, n184, n_249, n_290, n388, n412, n508, n538, n580, n686, n617, n_49, n_464, n_472, n_77, n_87, n658, n_123, n427, n_522, n_218, n_257, n_286, n_298, n_308, n_326, n_369, n_409, n551, n_544, n_483, n_532, n_584, n_596, n_19, n_499, n68, n241, n_268, n393, n513, n534, n576, n679, n685, n_173, n_230, n_272, n_315, n651, n_329, n_351, n432, n_422, n_459, n575, n_475, n_580, n168, n361, \ctoken_len[0], \ctoken_len[1], \ctoken_len[2], n_126, n_106, n_129, n407, n223, n_387, n489, n591, n_63, n_80, n_608, n_288, n_427, n_211, n_241, n365, n_363, n455, n495, n_486, n_508, n123, n182, n_339, n664, n_74, n_103, n_116, n_431, n_575, n_186, n_434, n_262, n_412, n_20, n468, n600, n_609, n638, n_70, n_305, n_494, n_238, n316, n_269, n_373, n_470, n_521, n389, n_43, n_449, n_189, n_332, n_280, n_90, n_120, n_278, n_348, n_385, n_452, n_497, n_513, n_67, n_50, n_113, n_382, n_275, n_517, n_398, n_393, n_243, n_150, n_164, n_224, n_304, n_509, n_552, n_235, n_380, n_198, n_35, n_40, n_144, n_340, n_418, n_448, n_482, n_572, n_549, n_354, n33, n_55, n_192, n_320, n_425, n_444, n_479, n_566, n_541, n_358, n_132, n_291, n_334, n_176, n_403, n_493, n_293, n_376, n_407, n_100, n_141, n_555, n_388, n_500, n_529, n_251, n_317, n_23;
	wire n33_key, n389_key, n316_key, n638_key, n600_key, n468_key, n317_key, n265_key, n275_key, n304_key, n345_key, n272_key, n307_key, n321_key, n262_key, n281_key, n328_key, n260_key, n274_key, n301_key, n311_key, n276_key, n323_key, n263_key, n314_key, n324_key, n331_key, n298_key, n346_key, n343_key, n337_key, n271_key, n279_key, n296_key, n284_key, n278_key, n312_key, n335_key, n302_key, n309_key, n289_key, n339_key, n350_key, n292_key, n258_key, n319_key, n341_key, n315_key, n270_key, n277_key, n318_key, n268_key, n330_key, n256_key, n269_key, n308_key, n347_key, n313_key, n273_key, n322_key, n326_key, n333_key, n288_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62;
	assign n_9 = ~\totalcoeffs[0];
	assign n28 = ( \totalcoeffs[0] & n_13 );
	assign n42 = ( \totalcoeffs[0] & \totalcoeffs[3] );
	assign n60 = ( \totalcoeffs[0] & n_22 );
	assign n75 = ( \totalcoeffs[0] & \trailingones[1] );
	assign n144 = ( \totalcoeffs[0] & \trailingones[0] );
	assign n172 = ( \totalcoeffs[0] & n171 );
	assign n195 = ( \totalcoeffs[0] & n194 );
	assign n202 = ( \totalcoeffs[0] & n201 );
	assign n203 = ( \totalcoeffs[0] & n_4 );
	assign n217 = ( \totalcoeffs[0] & \totalcoeffs[1] );
	assign n230 = ( \totalcoeffs[0] & n_179 );
	assign n317 = ( \totalcoeffs[0] & n_251 );
	assign n396 = ( \totalcoeffs[0] & n_323 );
	assign n441 = ( \totalcoeffs[0] & n_363 );
	assign n471 = ( \totalcoeffs[0] & n_389 );
	assign n480 = ( \totalcoeffs[0] & n170 );
	assign n522 = ( \totalcoeffs[0] & n_431 );
	assign n560 = ( \totalcoeffs[0] & n_464 );
	assign n643 = ( \totalcoeffs[0] & n_532 );
	assign n674 = ( \totalcoeffs[0] & n_561 );
	assign n_6 = ~\totalcoeffs[1];
	assign n25 = ( \totalcoeffs[1] & n_10 );
	assign n30 = ( \totalcoeffs[1] & n_13 );
	assign n37 = ( \totalcoeffs[1] & \totalcoeffs[2] );
	assign n45 = ( \totalcoeffs[1] & n_3 );
	assign n55 = ( \totalcoeffs[1] & n_43 );
	assign n56 = ( \totalcoeffs[1] & n_16 );
	assign n77 = ( \totalcoeffs[1] & n_60 );
	assign n105 = ( \totalcoeffs[1] & n_39 );
	assign n185 = ( \totalcoeffs[1] & n_144 );
	assign n206 = ( \totalcoeffs[1] & n_160 );
	assign n225 = ( \totalcoeffs[1] & \ctable[0] );
	assign n265 = ( \totalcoeffs[1] & n_211 );
	assign n275 = ( \totalcoeffs[1] & \trailingones[0] );
	assign n283 = ( \totalcoeffs[1] & n255 );
	assign n304 = ( \totalcoeffs[1] & n_241 );
	assign n320 = ( \totalcoeffs[1] & \trailingones[1] );
	assign n345 = ( \totalcoeffs[1] & n_280 );
	assign n371 = ( \totalcoeffs[1] & n_298 );
	assign n390 = ( \totalcoeffs[1] & n_317 );
	assign n414 = ( \totalcoeffs[1] & n290 );
	assign n501 = ( \totalcoeffs[1] & n_412 );
	assign n539 = ( \totalcoeffs[1] & n_448 );
	assign n577 = ( \totalcoeffs[1] & n_479 );
	assign n632 = ( \totalcoeffs[1] & n631 );
	assign n687 = ( \totalcoeffs[1] & n_572 );
	assign n_22 = ~\totalcoeffs[2];
	assign n62 = ( \totalcoeffs[2] & n_13 );
	assign n78 = ( \totalcoeffs[2] & n77 );
	assign n84 = ( n_6 & \totalcoeffs[2] );
	assign n95 = ( \totalcoeffs[2] & \trailingones[1] );
	assign n103 = ( \totalcoeffs[2] & n_3 );
	assign n158 = ( \totalcoeffs[2] & n_120 );
	assign n211 = ( \totalcoeffs[2] & n_165 );
	assign n243 = ( \totalcoeffs[2] & n_193 );
	assign n261 = ( \totalcoeffs[2] & n_4 );
	assign n272 = ( \totalcoeffs[2] & n_215 );
	assign n307 = ( \totalcoeffs[2] & n_243 );
	assign n321 = ( \totalcoeffs[2] & n320 );
	assign n325 = ( \totalcoeffs[2] & n125 );
	assign n353 = ( \totalcoeffs[2] & \ctable[1] );
	assign n366 = ( \totalcoeffs[2] & n_293 );
	assign n372 = ( \totalcoeffs[2] & n266 );
	assign n377 = ( \totalcoeffs[2] & n_305 );
	assign n399 = ( \totalcoeffs[2] & n398 );
	assign n436 = ( \totalcoeffs[2] & n_359 );
	assign n443 = ( \totalcoeffs[2] & n442 );
	assign n446 = ( \totalcoeffs[2] & n24 );
	assign n472 = ( \totalcoeffs[2] & n30 );
	assign n497 = ( \totalcoeffs[2] & n_236 );
	assign n506 = ( \totalcoeffs[2] & \trailingones[0] );
	assign n535 = ( \totalcoeffs[2] & n_444 );
	assign n578 = ( \totalcoeffs[2] & \totalcoeffs[3] );
	assign n593 = ( \totalcoeffs[2] & n_494 );
	assign n641 = ( \totalcoeffs[2] & n_530 );
	assign n645 = ( \totalcoeffs[2] & n_533 );
	assign n697 = ( \totalcoeffs[2] & n696 );
	assign n711 = ( \totalcoeffs[2] & n710 );
	assign n_3 = ~\totalcoeffs[3];
	assign n89 = ( \totalcoeffs[3] & n_70 );
	assign n110 = ( \totalcoeffs[3] & n_84 );
	assign n198 = ( \totalcoeffs[3] & \trailingones[0] );
	assign n214 = ( \totalcoeffs[3] & n213 );
	assign n226 = ( \totalcoeffs[3] & n_39 );
	assign n232 = ( \totalcoeffs[3] & n37 );
	assign n259 = ( \totalcoeffs[3] & n_205 );
	assign n262 = ( \totalcoeffs[3] & n_207 );
	assign n281 = ( \totalcoeffs[3] & n_224 );
	assign n310 = ( n_6 & \totalcoeffs[3] );
	assign n328 = ( \totalcoeffs[3] & n_262 );
	assign n352 = ( \totalcoeffs[3] & n_128 );
	assign n368 = ( \totalcoeffs[3] & n_294 );
	assign n386 = ( \totalcoeffs[3] & n_4 );
	assign n398 = ( \totalcoeffs[3] & n_54 );
	assign n413 = ( \totalcoeffs[3] & n_340 );
	assign n423 = ( \totalcoeffs[3] & n_99 );
	assign n490 = ( \totalcoeffs[3] & n_403 );
	assign n531 = ( \totalcoeffs[3] & n_372 );
	assign n545 = ( \totalcoeffs[3] & n_452 );
	assign n554 = ( n_22 & \totalcoeffs[3] );
	assign n568 = ( \totalcoeffs[3] & \ctable[0] );
	assign n571 = ( \totalcoeffs[3] & n491 );
	assign n677 = ( \totalcoeffs[3] & n_115 );
	assign n690 = ( \totalcoeffs[3] & n_575 );
	assign n_99 = ~\totalcoeffs[4];
	assign n127 = ( \totalcoeffs[4] & \trailingones[0] );
	assign n132 = ( \totalcoeffs[4] & \trailingones[1] );
	assign n293 = ( n_3 & \totalcoeffs[4] );
	assign n515 = ( n_6 & \totalcoeffs[4] );
	assign n603 = ( \totalcoeffs[4] & n_16 );
	assign n669 = ( \totalcoeffs[4] & n_558 );
	assign n691 = ( \totalcoeffs[4] & n_576 );
	assign n_4 = ~\ctable[0];
	assign n79 = ( \ctable[0] & n78 );
	assign n94 = ( \ctable[0] & n_74 );
	assign n130 = ( \ctable[0] & n_103 );
	assign n134 = ( \ctable[0] & \ctable[1] );
	assign n149 = ( \ctable[0] & n_113 );
	assign n162 = ( \ctable[0] & n_39 );
	assign n173 = ( n_9 & \ctable[0] );
	assign n192 = ( \ctable[0] & n146 );
	assign n231 = ( \ctable[0] & n_28 );
	assign n260 = ( \ctable[0] & n_206 );
	assign n274 = ( \ctable[0] & n_218 );
	assign n301 = ( \ctable[0] & n_238 );
	assign n311 = ( \ctable[0] & n_247 );
	assign n363 = ( \ctable[0] & \trailingones[0] );
	assign n367 = ( \ctable[0] & n_215 );
	assign n381 = ( \ctable[0] & \trailingones[1] );
	assign n439 = ( \ctable[0] & n320 );
	assign n448 = ( \ctable[0] & n_369 );
	assign n491 = ( n_22 & \ctable[0] );
	assign n561 = ( \ctable[0] & n_13 );
	assign n582 = ( \ctable[0] & n_483 );
	assign n610 = ( n_6 & \ctable[0] );
	assign n_54 = ~\ctable[1];
	assign n73 = ( \ctable[1] & n_57 );
	assign n91 = ( \ctable[1] & n_71 );
	assign n100 = ( \ctable[1] & n99 );
	assign n109 = ( n_22 & \ctable[1] );
	assign n128 = ( \ctable[1] & n127 );
	assign n131 = ( \ctable[1] & n_13 );
	assign n151 = ( \ctable[1] & \trailingones[1] );
	assign n170 = ( \ctable[1] & \trailingones[0] );
	assign n179 = ( n_9 & \ctable[1] );
	assign n210 = ( n_6 & \ctable[1] );
	assign n235 = ( \ctable[1] & n_183 );
	assign n266 = ( n_4 & \ctable[1] );
	assign n276 = ( \ctable[1] & n_219 );
	assign n282 = ( \ctable[1] & n_39 );
	assign n323 = ( \ctable[1] & n_257 );
	assign n329 = ( \ctable[1] & n_11 );
	assign n451 = ( \ctable[1] & n_373 );
	assign n499 = ( \ctable[1] & n_409 );
	assign n701 = ( \ctable[1] & n_585 );
	assign n_16 = ~\ctable[2];
	assign n51 = ( \ctable[2] & \trailingones[0] );
	assign n249 = ( \ctable[2] & n_198 );
	assign n457 = ( \ctable[2] & n_13 );
	assign n464 = ( \ctable[2] & n_382 );
	assign n675 = ( \ctable[2] & n_562 );
	assign n_39 = ~\trailingones[0];
	assign n81 = ( \trailingones[0] & n_63 );
	assign n102 = ( \trailingones[0] & n_80 );
	assign n150 = ( n_4 & \trailingones[0] );
	assign n154 = ( \trailingones[0] & n151 );
	assign n186 = ( n_54 & \trailingones[0] );
	assign n201 = ( n_22 & \trailingones[0] );
	assign n215 = ( n_9 & \trailingones[0] );
	assign n263 = ( \trailingones[0] & n_208 );
	assign n290 = ( \trailingones[0] & n_13 );
	assign n299 = ( \trailingones[0] & n75 );
	assign n314 = ( n_6 & \trailingones[0] );
	assign n324 = ( \trailingones[0] & n_258 );
	assign n331 = ( \trailingones[0] & n_264 );
	assign n356 = ( \trailingones[0] & \trailingones[1] );
	assign n445 = ( \trailingones[0] & n_366 );
	assign n458 = ( \trailingones[0] & n_377 );
	assign n520 = ( n_3 & \trailingones[0] );
	assign n564 = ( \trailingones[0] & n_467 );
	assign n586 = ( \trailingones[0] & n381 );
	assign n624 = ( \trailingones[0] & n_517 );
	assign n646 = ( \trailingones[0] & n_17 );
	assign n23 = ( n_6 & \trailingones[1] );
	assign n24 = ( n_9 & \trailingones[1] );
	assign n_13 = ~\trailingones[1];
	assign n41 = ( \trailingones[1] & n_28 );
	assign n53 = ( n_16 & \trailingones[1] );
	assign n161 = ( n_54 & \trailingones[1] );
	assign n174 = ( n_39 & \trailingones[1] );
	assign n238 = ( \trailingones[1] & n_186 );
	assign n255 = ( n_3 & \trailingones[1] );
	assign n401 = ( \trailingones[1] & n_326 );
	assign n452 = ( n_22 & \trailingones[1] );
	assign n484 = ( \trailingones[1] & n_398 );
	assign n525 = ( \trailingones[1] & n_434 );
	assign n636 = ( \trailingones[1] & n_525 );
	assign n36 = ( n_9 & n_24 );
	assign n63 = ( n_9 & n_6 );
	assign n70 = ( n_9 & n_22 );
	assign n74 = ( n_9 & n_13 );
	assign n98 = ( n_9 & n_3 );
	assign n107 = ( n_9 & n_83 );
	assign n116 = ( n_9 & n40 );
	assign n153 = ( n_9 & n_116 );
	assign n200 = ( n_9 & n_156 );
	assign n298 = ( n_9 & n_235 );
	assign n376 = ( n_9 & n_304 );
	assign n425 = ( n_9 & n227 );
	assign n442 = ( n_9 & n_333 );
	assign n461 = ( n_9 & n_380 );
	assign n474 = ( n_9 & n_54 );
	assign n485 = ( n_9 & n_39 );
	assign n543 = ( n_9 & n451 );
	assign n546 = ( n_9 & n146 );
	assign n562 = ( n_9 & n561 );
	assign n570 = ( n_9 & n_472 );
	assign n594 = ( n_9 & n593 );
	assign n609 = ( n_9 & n_505 );
	assign n654 = ( n_9 & n_544 );
	assign n142 = ( n_608 & n_9 & n_16 & n140 );
	assign n_14 = ~n28;
	assign n85 = ( n28 & n84 );
	assign n346 = ( n28 & n212 );
	assign n_30 = ~n42;
	assign n583 = ( n42 & n325 );
	assign n61 = ( n_47 & n60 );
	assign n596 = ( n60 & n595 );
	assign n_59 = ~n75;
	assign n343 = ( n51 & n75 );
	assign n145 = ( n95 & n144 );
	assign n462 = ( n144 & n320 );
	assign n_439 = ~n144;
	assign n_134 = ~n172;
	assign n_153 = ~n195;
	assign n_159 = ~n202;
	assign n_158 = ~n203;
	assign n337 = ( n203 & n_272 );
	assign n622 = ( n139 & n203 );
	assign n670 = ( n203 & n399 );
	assign n_169 = ~n217;
	assign n479 = ( n_39 & n217 );
	assign n_182 = ~n230;
	assign n_253 = ~n317_key;
	assign n418 = ~( n396 | n406 | n413 | n415 );
	assign n_364 = ~n441;
	assign n_390 = ~n471;
	assign n_394 = ~n480;
	assign n_437 = ~n522;
	assign n_465 = ~n560;
	assign n_537 = ~n643;
	assign n_619 = ~( n674 | n675 );
	assign n29 = ( n_6 & n_14 );
	assign n44 = ( n_6 & n_31 );
	assign n82 = ( n_6 & n_10 );
	assign n108 = ( n_6 & n_13 );
	assign n139 = ( n_6 & n_3 );
	assign n169 = ( n_6 & n_132 );
	assign n197 = ( n_6 & n_154 );
	assign n212 = ( n_6 & n_39 );
	assign n216 = ( n_6 & n_54 );
	assign n227 = ( n_6 & n_22 );
	assign n271 = ( n_6 & n_156 );
	assign n279 = ( n_6 & n174 );
	assign n362 = ( n_6 & n_291 );
	assign n406 = ( n_6 & n_332 );
	assign n435 = ( n_6 & n_4 );
	assign n509 = ( n_6 & n_418 );
	assign n553 = ( n_6 & n_459 );
	assign n585 = ( n_6 & n_486 );
	assign n640 = ( n_6 & n_236 );
	assign n659 = ( n_6 & n_549 );
	assign n699 = ( n_6 & n_584 );
	assign n296 = ( n_612 & n_22 & n_6 & n293 );
	assign n_12 = ~n25;
	assign n_17 = ~n30;
	assign n96 = ( n_22 & n30 );
	assign n247 = ( n30 & n201 );
	assign n487 = ( n30 & n486 );
	assign n_26 = ~n37;
	assign n627 = ( n37 & n626 );
	assign n_33 = ~n45;
	assign n_45 = ~n55;
	assign n_44 = ~n56;
	assign n92 = ( n40 & n77 );
	assign n_82 = ~n105;
	assign n_145 = ~n185;
	assign n_162 = ~n206;
	assign n_177 = ~n225;
	assign n_212 = ~n265_key;
	assign n_219 = ~n275_key;
	assign n284 = ( n282 & n283 );
	assign n_503 = ~n283;
	assign n_244 = ~n304_key;
	assign n_265 = ~n320;
	assign n660 = ( n320 & n546 );
	assign n_281 = ~n345_key;
	assign n_299 = ~n371;
	assign n_321 = ~n390;
	assign n415 = ( n266 & n414 );
	assign n_419 = ~n501;
	assign n_462 = ~n539;
	assign n_489 = ~n577;
	assign n_523 = ~n632;
	assign n_620 = ~( n687 | n699 );
	assign n34 = ( n_22 & n_23 );
	assign n35 = ( n_22 & n_4 );
	assign n40 = ( n_22 & n_3 );
	assign n90 = ( n_22 & n_14 );
	assign n140 = ( n_22 & n139 );
	assign n146 = ( n_22 & n_39 );
	assign n177 = ( n_22 & n_136 );
	assign n180 = ( n_22 & n_137 );
	assign n199 = ( n_22 & n_155 );
	assign n278 = ( n_22 & n_221 );
	assign n312 = ( n_22 & n125 );
	assign n335 = ( n_22 & n_269 );
	assign n359 = ( n_22 & n293 );
	assign n378 = ( n_22 & n363 );
	assign n384 = ( n_22 & n_310 );
	assign n408 = ( n_22 & n_334 );
	assign n465 = ( n_22 & n464 );
	assign n482 = ( n_22 & n_395 );
	assign n505 = ( n_22 & n504 );
	assign n529 = ( n_22 & n_438 );
	assign n542 = ( n_22 & n541 );
	assign n579 = ( n_22 & n_30 );
	assign n621 = ( n_22 & n620 );
	assign n680 = ( n_22 & n_566 );
	assign n694 = ( n_22 & n_580 );
	assign n220 = ( n_610 & n_22 & n_170 & n_169 );
	assign n614 = ( n_22 & n_508 & n_242 & n_203 );
	assign n64 = ( n62 & n63 );
	assign n187 = ( n62 & n186 );
	assign n_258 = ~n62;
	assign n459 = ( n84 & n_378 );
	assign n_75 = ~n95;
	assign n302 = ( n_4 & n95 );
	assign n565 = ( n95 & n162 );
	assign n657 = ( n95 & n485 );
	assign n104 = ( n23 & n103 );
	assign n616 = ( n103 & n_509 );
	assign n_562 = ~n103;
	assign n_122 = ~n158;
	assign n_166 = ~n211;
	assign n_194 = ~n243;
	assign n422 = ( n_99 & n243 );
	assign n_207 = ~n261;
	assign n_217 = ~n272_key;
	assign n_245 = ~n307_key;
	assign n_256 = ~n321_key;
	assign n_260 = ~n325;
	assign n_285 = ~n353;
	assign n_297 = ~n366;
	assign n_300 = ~n372;
	assign n_306 = ~n377;
	assign n_325 = ~n399;
	assign n681 = ( n_372 & n399 );
	assign n_360 = ~n436;
	assign n_365 = ~n443;
	assign n_368 = ~n446;
	assign n_391 = ~n472;
	assign n_408 = ~n497;
	assign n550 = ( n497 & n_455 );
	assign n507 = ( n24 & n506 );
	assign n_543 = ~n506;
	assign n_445 = ~n535;
	assign n_481 = ~n578;
	assign n587 = ( n578 & n586 );
	assign n_531 = ~n641;
	assign n_535 = ~n645;
	assign n_583 = ~n697;
	assign n_595 = ~n711;
	assign n22 = ( n_3 & n_4 );
	assign n67 = ( n_3 & n_50 );
	assign n191 = ( n_3 & n_150 );
	assign n193 = ( n_3 & n_39 );
	assign n309 = ( n_3 & n_246 );
	assign n383 = ( n_3 & n_309 );
	assign n391 = ( n_3 & n266 );
	assign n469 = ( n_3 & n_388 );
	assign n530 = ( n_3 & n356 );
	assign n536 = ( n_3 & n126 );
	assign n567 = ( n_3 & n_470 );
	assign n676 = ( n_3 & n_333 );
	assign n684 = ( n_3 & n_568 );
	assign n692 = ( n_3 & n_577 );
	assign n121 = ~( n89 | n102 | n115 | n118 );
	assign n_85 = ~n110;
	assign n_155 = ~n198;
	assign n_171 = ~n214;
	assign n228 = ( n226 & n227 );
	assign n_311 = ~n226;
	assign n_181 = ~n232;
	assign n236 = ( n162 & n232 );
	assign n_206 = ~n259;
	assign n_208 = ~n262_key;
	assign n_614 = ~n281_key;
	assign n_247 = ~n310;
	assign n633 = ( n_157 & n310 );
	assign n_270 = ~n328_key;
	assign n_284 = ~n352;
	assign n_296 = ~n368;
	assign n_313 = ~n386;
	assign n650 = ( n386 & n_538 );
	assign n_327 = ~n398;
	assign n523 = ( n215 & n398 );
	assign n_350 = ~n423;
	assign n431 = ( n423 & n_355 );
	assign n710 = ( n423 & n_594 );
	assign n_421 = ~n490;
	assign n_440 = ~n531;
	assign n_458 = ~n545;
	assign n556 = ( n554 & n555 );
	assign n574 = ( n554 & n561 );
	assign n_471 = ~n568;
	assign n_474 = ~n571;
	assign n_563 = ~n677;
	assign n_578 = ~n690;
	assign n124 = ( n_99 & n_100 );
	assign n160 = ( n_99 & n_123 );
	assign n189 = ( n_99 & n_147 );
	assign n240 = ( n_99 & n_189 );
	assign n289 = ( n_99 & n_230 );
	assign n339 = ( n_99 & n_275 );
	assign n355 = ( n_99 & n_286 );
	assign n374 = ( n_99 & n_301 );
	assign n419 = ( n_99 & n_345 );
	assign n514 = ( n_99 & n_425 );
	assign n601 = ( n_99 & n_500 );
	assign n665 = ( n_99 & n_555 );
	assign n253 = ( n_609 & n22 & n_54 & n_99 );
	assign n350 = ( n_611 & n342 & n40 & n_99 );
	assign n_124 = ~n127;
	assign n_105 = ~n132;
	assign n_349 = ~n293;
	assign n516 = ( n116 & n515 );
	assign n666 = ( n22 & n603 );
	assign n605 = ( n35 & n98 & n216 & n603 );
	assign n_618 = ~( n669 | n672 );
	assign n_577 = ~n691;
	assign n52 = ( n_4 & n51 );
	assign n57 = ( n_4 & n_13 );
	assign n72 = ( n_4 & n_56 );
	assign n87 = ( n_4 & n_67 );
	assign n115 = ( n_4 & n_90 );
	assign n222 = ( n_4 & n_173 );
	assign n292 = ( n_4 & n291 );
	assign n342 = ( n_4 & n_54 );
	assign n478 = ( n_4 & n_393 );
	assign n559 = ( n_4 & n_463 );
	assign n625 = ( n_4 & n_170 );
	assign n682 = ( n_4 & n681 );
	assign n700 = ( n_4 & n_562 );
	assign n_62 = ~n79;
	assign n_78 = ~n94;
	assign n_108 = ~n130;
	assign n_107 = ~n134;
	assign \coeff_token[4] = ( n134 & n428 );
	assign \coeff_token[5] = ( n134 & n433 );
	assign n_121 = ~n149;
	assign n_125 = ~n162;
	assign n175 = ( n173 & n174 );
	assign n_157 = ~n173;
	assign n_152 = ~n192;
	assign n392 = ( n192 & n216 );
	assign n_180 = ~n231;
	assign n_209 = ~n260_key;
	assign n_613 = ~n274_key;
	assign n_239 = ~n301_key;
	assign n_248 = ~n311_key;
	assign n364 = ( n161 & n363 );
	assign n_336 = ~n363;
	assign n_294 = ~n367;
	assign n382 = ( n_39 & n381 );
	assign n_335 = ~n381;
	assign n_362 = ~n439;
	assign n_371 = ~n448;
	assign n492 = ( n_60 & n491 );
	assign n607 = ( n227 & n561 );
	assign n_484 = ~n582;
	assign n_507 = ~n610;
	assign n69 = ( n_54 & n_55 );
	assign n126 = ( n_54 & n125 );
	assign n164 = ( n_54 & n_126 );
	assign n178 = ( n_54 & n_39 );
	assign n209 = ( n_54 & n_164 );
	assign n258 = ( n_54 & n257 );
	assign n319 = ( n_54 & n_254 );
	assign n385 = ( n_54 & n_311 );
	assign n409 = ( n_54 & n_335 );
	assign n438 = ( n_54 & n437 );
	assign n493 = ( n_54 & n_207 );
	assign n533 = ( n_54 & n_441 );
	assign n541 = ( n_54 & n_449 );
	assign n549 = ( n_54 & n_151 );
	assign n590 = ( n_54 & n_490 );
	assign n639 = ( n_54 & n_529 );
	assign n644 = ( n_54 & n_82 );
	assign n663 = ( n_54 & n662 );
	assign n683 = ( n_54 & n_567 );
	assign n_61 = ~n73;
	assign n_72 = ~n91;
	assign n_79 = ~n100;
	assign n_84 = ~n109;
	assign n_102 = ~n128;
	assign n_104 = ~n131;
	assign n_115 = ~n151;
	assign n_133 = ~n170;
	assign n526 = ( n_13 & n170 );
	assign n_137 = ~n179;
	assign n_165 = ~n210;
	assign n_184 = ~n235;
	assign n267 = ( n_39 & n266 );
	assign n397 = ( n_28 & n266 );
	assign n402 = ( n_13 & n266 );
	assign n_220 = ~n276_key;
	assign n_432 = ~n282;
	assign n555 = ( n_13 & n282 );
	assign n_261 = ~n323_key;
	assign n_263 = ~n329;
	assign n647 = ( n329 & n_534 );
	assign n454 = ( n451 & n453 );
	assign n_411 = ~n499;
	assign n_617 = ~n701;
	assign n31 = ( n_16 & n_17 );
	assign n48 = ( n_16 & n_35 );
	assign n122 = ( n_16 & n_95 );
	assign n242 = ( n_16 & n_192 );
	assign n341 = ( n_16 & n_278 );
	assign \coeff_token[3] = ( n_16 & n_348 );
	assign n428 = ( n_16 & n_354 );
	assign n433 = ( n_16 & n_358 );
	assign n456 = ( n_16 & n_376 );
	assign n512 = ( n_16 & n_422 );
	assign n518 = ( n_16 & n_427 );
	assign n592 = ( n_16 & n_493 );
	assign n652 = ( n_16 & n_541 );
	assign n671 = ( n_16 & n_559 );
	assign n673 = ( n_16 & n_558 );
	assign n713 = ( n_16 & n_596 );
	assign n595 = ( n_13 & n51 );
	assign n_200 = ~n249;
	assign n_377 = ~n457;
	assign n50 = ( n_39 & n_40 );
	assign n83 = ( n_39 & n_64 );
	assign n113 = ( n_39 & n_87 );
	assign n117 = ( n_39 & n108 );
	assign n125 = ( n_39 & n_13 );
	assign n136 = ( n_39 & n135 );
	assign n155 = ( n_39 & n57 );
	assign n246 = ( n_39 & n245 );
	assign n404 = ( n_39 & n_329 );
	assign n496 = ( n_39 & n_407 );
	assign n502 = ( n_39 & n_413 );
	assign n573 = ( n_39 & n_475 );
	assign n619 = ( n_39 & n_513 );
	assign n695 = ( n_39 & n_335 );
	assign n708 = ( n_39 & n_18 );
	assign n_68 = ~n81;
	assign n_114 = ~n150;
	assign n181 = ( n150 & n_138 );
	assign n_117 = ~n154;
	assign n_215 = ~n186;
	assign n_205 = ~n201;
	assign n634 = ( n201 & n633 );
	assign n_170 = ~n215;
	assign n678 = ( n215 & n_563 );
	assign n688 = ( n215 & n_573 );
	assign n_210 = ~n263_key;
	assign n_231 = ~n290;
	assign n_237 = ~n299;
	assign n315 = ( n41 & n314_key );
	assign n_255 = ~n314_key;
	assign n_259 = ~n324_key;
	assign n_267 = ~n331_key;
	assign n357 = ( n342 & n356 );
	assign n_372 = ~n356;
	assign n_370 = ~n445;
	assign n_378 = ~n458;
	assign n_430 = ~n520;
	assign n_468 = ~n564;
	assign n_567 = ~n586;
	assign n_519 = ~n624;
	assign n_534 = ~n646;
	assign n_11 = ~n23;
	assign n71 = ( n23 & n70 );
	assign n_10 = ~n24;
	assign n494 = ( n24 & n_404 );
	assign n39 = ( n_13 & n_27 );
	assign n183 = ( n_13 & n_141 );
	assign n224 = ( n_13 & n_176 );
	assign n270 = ( n_13 & n_214 );
	assign n277 = ( n_13 & n_220 );
	assign n380 = ( n_13 & n_308 );
	assign n394 = ( n_13 & n_320 );
	assign n437 = ( n_13 & n_360 );
	assign n504 = ( n_13 & n_415 );
	assign n548 = ( n_13 & n_454 );
	assign n629 = ( n_13 & n_521 );
	assign n656 = ( n_13 & n_546 );
	assign n_29 = ~n41;
	assign n_42 = ~n53;
	assign n_128 = ~n161;
	assign n_202 = ~n174;
	assign n_188 = ~n238;
	assign n_203 = ~n255;
	assign n_330 = ~n401;
	assign n_374 = ~n452;
	assign n_400 = ~n484;
	assign n_435 = ~n525;
	assign n_527 = ~n636;
	assign n_25 = ~n36;
	assign n_193 = ~n63;
	assign n430 = ( n63 & n359 );
	assign n167 = ( n70 & n166 );
	assign n_58 = ~n74;
	assign n147 = ( n74 & n146 );
	assign n99 = ( n_77 & n98 );
	assign n_514 = ~n98;
	assign n_88 = ~n107;
	assign n118 = ( n116 & n117 );
	assign n_119 = ~n153;
	assign n_161 = ~n200;
	assign n_276 = ~n298_key;
	assign n_346 = ~n376;
	assign n426 = ( n_351 & n425 );
	assign n_355 = ~n425;
	assign n667 = ( n425 & n666 );
	assign n_383 = ~n461;
	assign n476 = ( n474 & n475 );
	assign n_413 = ~n474;
	assign n_399 = ~n485;
	assign n_451 = ~n543;
	assign n_453 = ~n546;
	assign n_466 = ~n562;
	assign n_473 = ~n570;
	assign n_495 = ~n594;
	assign n_512 = ~n609;
	assign n_545 = ~n654;
	assign \coeff_token[0] = ( n124 | n142 );
	assign n_66 = ~n85;
	assign n_282 = ~n346_key;
	assign n43 = ( n_29 & n_30 );
	assign n_485 = ~n583;
	assign n_48 = ~n61;
	assign n_496 = ~n596;
	assign n76 = ( n_58 & n_59 );
	assign n_279 = ~n343_key;
	assign n_111 = ~n145;
	assign n_381 = ~n462;
	assign n532 = ( n_439 & n_440 );
	assign n176 = ( n_134 & n_135 );
	assign n196 = ( n_152 & n_153 );
	assign n205 = ( n_159 & n204 );
	assign n655 = ( n_159 & n_545 );
	assign n204 = ( n_157 & n_158 );
	assign n486 = ( n_158 & n_399 );
	assign n503 = ( n_158 & n_414 );
	assign n_274 = ~n337_key;
	assign n_516 = ~n622;
	assign n_559 = ~n670;
	assign n244 = ( n90 & n_169 );
	assign n_396 = ~n479;
	assign n234 = ( n_182 & n233 );
	assign n318 = ( n_252 & n_253 );
	assign n_345 = ~n418;
	assign n444 = ( n_364 & n_365 );
	assign n473 = ( n_390 & n_391 );
	assign n481 = ( n_82 & n_394 );
	assign n547 = ( n_394 & n_453 );
	assign n528 = ( n_437 & n527 );
	assign n563 = ( n_465 & n_466 );
	assign n649 = ( n_537 & n648 );
	assign \ctoken_len[3] = ( n_617 & n_618 & n_619 & n_620 );
	assign n_18 = ~n29;
	assign n_32 = ~n44;
	assign n_64 = ~n82;
	assign n111 = ( n108 & n_85 );
	assign n_242 = ~n108;
	assign n268 = ( n139 & n267 );
	assign n_148 = ~n169;
	assign n_163 = ~n197;
	assign n_167 = ~n212;
	assign n598 = ( n216 & n_497 );
	assign n_610 = ~n216;
	assign n_216 = ~n271_key;
	assign n_223 = ~n279_key;
	assign n_302 = ~n362;
	assign n_359 = ~n435;
	assign n_420 = ~n509;
	assign n_460 = ~n553;
	assign n_487 = ~n585;
	assign n_530 = ~n640;
	assign n_550 = ~n659;
	assign n_234 = ~n296_key;
	assign n26 = ( n_11 & n_12 );
	assign n709 = ( n_12 & n_593 );
	assign n330 = ( n_17 & n_263 );
	assign n_76 = ~n96;
	assign n_197 = ~n247;
	assign n_401 = ~n487;
	assign n38 = ( n_25 & n_26 );
	assign n_520 = ~n627;
	assign n46 = ( n_32 & n_33 );
	assign n256 = ( n_33 & n_202 );
	assign n59 = ( n_45 & n_46 );
	assign n58 = ( n_44 & n57 );
	assign n_73 = ~n92;
	assign n106 = ( n_81 & n_82 );
	assign n188 = ( n_145 & n_146 );
	assign n207 = ( n_161 & n_162 );
	assign n229 = ( n_177 & n_178 );
	assign n269 = ( n_212 & n_213 );
	assign n_615 = ~n284_key;
	assign n608 = ( n_503 & n_504 );
	assign n308 = ( n_244 & n_245 );
	assign n332 = ( n_242 & n_265 );
	assign n410 = ( n_265 & n_336 );
	assign n470 = ( n_367 & n_265 );
	assign n_551 = ~n660;
	assign n347 = ( n_281 & n_282 );
	assign n373 = ( n_299 & n_300 );
	assign n395 = ( n_321 & n_322 );
	assign n510 = ( n_419 & n_420 );
	assign n558 = ( n_462 & n557 );
	assign n589 = ( n_489 & n588 );
	assign n635 = ( n_523 & n_524 );
	assign n_36 = ~n34;
	assign n_24 = ~n35;
	assign n_28 = ~n40;
	assign n_71 = ~n90;
	assign n_558 = ~n140;
	assign n_542 = ~n146;
	assign n_142 = ~n177;
	assign n_138 = ~n180;
	assign n_156 = ~n199;
	assign n_222 = ~n278_key;
	assign n313 = ( n_248 & n312_key );
	assign n_271 = ~n335_key;
	assign n360 = ( n_288 & n359 );
	assign n_307 = ~n378;
	assign n_314 = ~n384;
	assign n_338 = ~n408;
	assign n_384 = ~n465;
	assign n_397 = ~n482;
	assign n_416 = ~n505;
	assign n_447 = ~n529;
	assign n_450 = ~n542;
	assign n_480 = ~n579;
	assign n_515 = ~n621;
	assign n_571 = ~n680;
	assign n_582 = ~n694;
	assign n_172 = ~n220;
	assign n_510 = ~n614;
	assign n65 = ( n52 & n64 );
	assign n_199 = ~n64;
	assign n_146 = ~n187;
	assign n453 = ( n_258 & n_374 );
	assign n569 = ( n_258 & n_471 );
	assign n_379 = ~n459;
	assign n97 = ( n_75 & n_76 );
	assign n112 = ( n_75 & n_86 );
	assign n_240 = ~n302_key;
	assign n_469 = ~n565;
	assign n_548 = ~n657;
	assign n_81 = ~n104;
	assign n_511 = ~n616;
	assign n159 = ( n_121 & n_122 );
	assign n213 = ( n_166 & n_167 );
	assign n245 = ( n_194 & n_195 );
	assign n_352 = ~n422;
	assign n630 = ( n_207 & n_471 );
	assign n273 = ( n_216 & n_217 );
	assign n322 = ( n_255 & n_256 );
	assign n326 = ( n_259 & n_260 );
	assign n354 = ( n_284 & n_285 );
	assign n370 = ( n_297 & n369 );
	assign n379 = ( n_306 & n_307 );
	assign n400 = ( n_324 & n_325 );
	assign n447 = ( n_367 & n_368 );
	assign n498 = ( n_237 & n_408 );
	assign n_457 = ~n550;
	assign n_417 = ~n507;
	assign n653 = ( n_542 & n_543 );
	assign n537 = ( n_445 & n_446 );
	assign n581 = ( n_481 & n_482 );
	assign n_488 = ~n587;
	assign n642 = ( n_263 & n_531 );
	assign n648 = ( n_535 & n_536 );
	assign n698 = ( n_582 & n_583 );
	assign n712 = ( n_356 & n_595 );
	assign n27 = ( n22 & n26 );
	assign n599 = ( n22 & n598 );
	assign n_506 = ~n22;
	assign n662 = ( n22 & n_552 );
	assign n_52 = ~n67;
	assign n_190 = ~n191;
	assign n_151 = ~n193;
	assign n333 = ( n193 & n_266 );
	assign n_252 = ~n309_key;
	assign n_310 = ~n383;
	assign n_318 = ~n391;
	assign n_423 = ~n469;
	assign n_442 = ~n530;
	assign n_446 = ~n536;
	assign n_478 = ~n567;
	assign n_564 = ~n676;
	assign n696 = ( n676 & n_581 );
	assign n_570 = ~n684;
	assign n_579 = ~n692;
	assign n_95 = ~n121;
	assign n221 = ( n_171 & n_172 );
	assign n_178 = ~n228;
	assign n233 = ( n_180 & n_181 );
	assign n_185 = ~n236;
	assign n631 = ( n_206 & n_522 );
	assign n288 = ( n_613 & n_614 & n_615 & n_616 );
	assign n336 = ( n_270 & n_271 );
	assign n369 = ( n_295 & n_296 );
	assign n387 = ( n_312 & n_313 );
	assign n_540 = ~n650;
	assign n403 = ( n_327 & n_328 );
	assign n_433 = ~n523;
	assign n424 = ( n_349 & n_350 );
	assign n_357 = ~n431;
	assign n511 = ( n_421 & n510 );
	assign n552 = ( n_458 & n551 );
	assign n_461 = ~n556;
	assign n_477 = ~n574;
	assign n626 = ( n_471 & n_518 );
	assign n572 = ( n_473 & n_474 );
	assign n693 = ( n_578 & n_579 );
	assign n_130 = ~n160;
	assign n_149 = ~n189;
	assign n_191 = ~n240;
	assign n_233 = ~n289_key;
	assign n_277 = ~n339_key;
	assign n_289 = ~n355;
	assign n_303 = ~n374;
	assign n_347 = ~n419;
	assign n_428 = ~n514;
	assign n_501 = ~n601;
	assign n_556 = ~n665;
	assign \coeff_token[1] = ( n242 | n253 );
	assign \coeff_token[2] = ( n341_key | n350_key );
	assign n163 = ( n_124 & n_125 );
	assign n133 = ( n_104 & n_105 );
	assign n165 = ( n_105 & n_127 );
	assign n_426 = ~n516;
	assign n_502 = ~n605;
	assign n_41 = ~n52;
	assign n_333 = ~n57;
	assign n_57 = ~n72;
	assign n_69 = ~n87;
	assign n_175 = ~n222;
	assign n_612 = ~n292_key;
	assign n467 = ( n342 & n_385 );
	assign n_576 = ~n342;
	assign \ctoken_len[4] = ( n342 & n713 );
	assign n_402 = ~n478;
	assign n_491 = ~n559;
	assign n_518 = ~n625;
	assign n_569 = ~n682;
	assign n_585 = ~n700;
	assign n80 = ( n_61 & n_62 );
	assign n101 = ( n_78 & n_79 );
	assign n137 = ( n_108 & n_109 );
	assign n135 = ( n_106 & n_107 );
	assign n358 = ( n_107 & n_287 );
	assign n517 = ( n_107 & n_426 );
	assign n_135 = ~n175;
	assign n_319 = ~n392;
	assign n264 = ( n_209 & n_210 );
	assign n303 = ( n_239 & n_240 );
	assign n_292 = ~n364;
	assign n_309 = ~n382;
	assign n440 = ( n_361 & n_362 );
	assign n449 = ( n_370 & n_371 );
	assign n_405 = ~n492;
	assign n_504 = ~n607;
	assign n584 = ( n_484 & n_485 );
	assign n611 = ( n_506 & n_507 );
	assign n_96 = ~n69;
	assign n_101 = ~n126;
	assign n_127 = ~n164;
	assign n_139 = ~n178;
	assign n_174 = ~n209;
	assign n_616 = ~( n258_key | n270_key );
	assign n_273 = ~n319_key;
	assign n_312 = ~n385;
	assign n411 = ( n409 & n_337 );
	assign n_573 = ~n409;
	assign n_361 = ~n438;
	assign n_404 = ~n493;
	assign n_443 = ~n533;
	assign n_455 = ~n549;
	assign n_492 = ~n590;
	assign n_539 = ~n639;
	assign n_533 = ~n644;
	assign n_554 = ~n663;
	assign n_568 = ~n683;
	assign n93 = ( n_72 & n_73 );
	assign n129 = ( n_101 & n_102 );
	assign n152 = ( n_114 & n_115 );
	assign n521 = ( n_115 & n_430 );
	assign n689 = ( n_115 & n_574 );
	assign n171 = ( n_116 & n_133 );
	assign n_436 = ~n526;
	assign n237 = ( n_184 & n_185 );
	assign n_295 = ~n267;
	assign n_324 = ~n397;
	assign n_328 = ~n402;
	assign n524 = ( n_432 & n_433 );
	assign n327 = ( n_261 & n326_key );
	assign n_536 = ~n647;
	assign n_375 = ~n454;
	assign n500 = ( n_410 & n_411 );
	assign n32 = ( n_18 & n31 );
	assign n_37 = ~n48;
	assign n_97 = ~n122;
	assign n_386 = ~n456;
	assign n_424 = ~n512;
	assign n_429 = ~n518;
	assign n_498 = ~n592;
	assign n_553 = ~n652;
	assign n_560 = ~n671;
	assign n_561 = ~n673;
	assign n250 = ( n_199 & n_200 );
	assign n_51 = ~n50;
	assign n_65 = ~n83;
	assign n_89 = ~n113;
	assign n_367 = ~n117;
	assign n_236 = ~n125;
	assign n_109 = ~n136;
	assign n_118 = ~n155;
	assign n_196 = ~n246;
	assign n_331 = ~n404;
	assign n_410 = ~n496;
	assign n_414 = ~n502;
	assign n_476 = ~n573;
	assign n_528 = ~n619;
	assign n_581 = ~n695;
	assign n_593 = ~n708;
	assign n88 = ( n_68 & n_69 );
	assign n194 = ( n_114 & n_151 );
	assign n_140 = ~n181;
	assign n156 = ( n_117 & n_118 );
	assign n_524 = ~n634;
	assign n_565 = ~n678;
	assign n_574 = ~n688;
	assign n291 = ( n_139 & n_231 );
	assign n305 = ( n_202 & n_231 );
	assign n300 = ( n_236 & n_237 );
	assign n_250 = ~n315_key;
	assign n334 = ( n_267 & n_268 );
	assign n_287 = ~n357;
	assign n450 = ( n_236 & n_372 );
	assign n566 = ( n_468 & n_469 );
	assign n628 = ( n_519 & n_520 );
	assign n_56 = ~n71;
	assign n_406 = ~n494;
	assign n_34 = ~n39;
	assign n_143 = ~n183;
	assign n_187 = ~n224;
	assign n_221 = ~n277_key;
	assign n_316 = ~n380;
	assign n_322 = ~n394;
	assign n_456 = ~n548;
	assign n_526 = ~n629;
	assign n_547 = ~n656;
	assign n54 = ( n_41 & n_42 );
	assign n166 = ( n_128 & n_129 );
	assign n540 = ( n_58 & n_202 );
	assign n239 = ( n_187 & n_188 );
	assign n257 = ( n_203 & n_204 );
	assign n405 = ( n_330 & n_331 );
	assign n488 = ( n_400 & n_401 );
	assign n527 = ( n_435 & n_436 );
	assign n637 = ( n_526 & n_527 );
	assign n_356 = ~n430;
	assign n_131 = ~n167;
	assign n344 = ( n_58 & n_279 );
	assign n_112 = ~n147;
	assign n620 = ( n_514 & n_508 );
	assign n114 = ( n_88 & n_89 );
	assign n157 = ( n_119 & n156 );
	assign n340 = ( n_276 & n_277 );
	assign n420 = ( n_346 & n_347 );
	assign n_353 = ~n426;
	assign n_557 = ~n667;
	assign n466 = ( n_383 & n_384 );
	assign n_392 = ~n476;
	assign n544 = ( n_450 & n_451 );
	assign n597 = ( n_495 & n_496 );
	assign n618 = ( n_512 & n617 );
	assign n86 = ( n_65 & n_66 );
	assign n_31 = ~n43;
	assign n66 = ( n_48 & n_49 );
	assign n_60 = ~n76;
	assign n148 = ( n_111 & n_112 );
	assign n463 = ( n_236 & n_381 );
	assign n_441 = ~n532;
	assign n_136 = ~n176;
	assign n_154 = ~n196;
	assign n_160 = ~n205;
	assign n_546 = ~n655;
	assign n_415 = ~n503;
	assign n338 = ( n_273 & n_274 );
	assign n623 = ( n_515 & n_516 );
	assign n_195 = ~n244;
	assign n483 = ( n_396 & n_397 );
	assign n_183 = ~n234;
	assign n_254 = ~n318_key;
	assign n_366 = ~n444;
	assign n477 = ( n473 & n_392 );
	assign n_395 = ~n481;
	assign n_454 = ~n547;
	assign n_438 = ~n528;
	assign n_467 = ~n563;
	assign n_538 = ~n649;
	assign n_86 = ~n111;
	assign n306 = ( n_242 & n305 );
	assign n_213 = ~n268_key;
	assign n190 = ( n_148 & n_149 );
	assign n208 = ( n_163 & n207 );
	assign n475 = ( n_167 & n332 );
	assign n280 = ( n_222 & n_223 );
	assign n375 = ( n_302 & n_303 );
	assign n615 = ( n332 & n_359 );
	assign n557 = ( n_460 & n_461 );
	assign n588 = ( n_487 & n_488 );
	assign n672 = ( n_530 & n_560 );
	assign n661 = ( n_550 & n_551 );
	assign n297 = ( n_233 & n_234 );
	assign n_594 = ~n709;
	assign n_264 = ~n330_key;
	assign n460 = ( n_76 & n_379 );
	assign n248 = ( n_196 & n_197 );
	assign n_27 = ~n38;
	assign n47 = ( n_34 & n46 );
	assign n_204 = ~n256_key;
	assign n_47 = ~n59;
	assign n_46 = ~n58;
	assign n_83 = ~n106;
	assign n_147 = ~n188;
	assign n_179 = ~n229;
	assign n_214 = ~n269_key;
	assign n_505 = ~n608;
	assign n_246 = ~n308_key;
	assign n_266 = ~n332;
	assign n_337 = ~n410;
	assign n_389 = ~n470;
	assign n_611 = ~n347_key;
	assign n_301 = ~n373;
	assign n_323 = ~n395;
	assign n_463 = ~n558;
	assign n_490 = ~n589;
	assign n_525 = ~n635;
	assign n49 = ( n_36 & n_37 );
	assign n184 = ( n_142 & n_143 );
	assign n_249 = ~n313_key;
	assign n_290 = ~n360;
	assign n388 = ( n_314 & n_315 );
	assign n412 = ( n_338 & n_339 );
	assign n508 = ( n_416 & n_417 );
	assign n538 = ( n_447 & n537 );
	assign n580 = ( n_373 & n_480 );
	assign n686 = ( n_571 & n685 );
	assign n617 = ( n_510 & n_511 );
	assign n_49 = ~n65;
	assign n_464 = ~n453;
	assign n_472 = ~n569;
	assign n_77 = ~n97;
	assign n_87 = ~n112;
	assign n658 = ( n_547 & n_548 );
	assign n_123 = ~n159;
	assign n427 = ( n_352 & n_353 );
	assign n_522 = ~n630;
	assign n_218 = ~n273_key;
	assign n_257 = ~n322_key;
	assign n_286 = ~n354;
	assign n_298 = ~n370;
	assign n_308 = ~n379;
	assign n_326 = ~n400;
	assign n_369 = ~n447;
	assign n_409 = ~n498;
	assign n551 = ( n_456 & n_457 );
	assign n_544 = ~n653;
	assign n_483 = ~n581;
	assign n_532 = ~n642;
	assign n_584 = ~n698;
	assign n_596 = ~n712;
	assign n_19 = ~n27;
	assign n_499 = ~n599;
	assign n68 = ( n_51 & n_52 );
	assign n241 = ( n_190 & n_191 );
	assign n_268 = ~n333_key;
	assign n393 = ( n_318 & n_319 );
	assign n513 = ( n_423 & n_424 );
	assign n534 = ( n_442 & n_443 );
	assign n576 = ( n_478 & n575 );
	assign n679 = ( n_564 & n_565 );
	assign n685 = ( n_569 & n_570 );
	assign n_173 = ~n221;
	assign n_230 = ~n288_key;
	assign n_272 = ~n336;
	assign n_315 = ~n387;
	assign n651 = ( n_539 & n_540 );
	assign n_329 = ~n403;
	assign n_351 = ~n424;
	assign n432 = ( n_356 & n_357 );
	assign n_422 = ~n511;
	assign n_459 = ~n552;
	assign n575 = ( n_476 & n_477 );
	assign n_475 = ~n572;
	assign n_580 = ~n693;
	assign n168 = ( n_130 & n_131 );
	assign n361 = ( n_289 & n_290 );
	assign \ctoken_len[0] = ( n_428 & n_429 );
	assign \ctoken_len[1] = ( n_501 & n_502 );
	assign \ctoken_len[2] = ( n_556 & n_557 );
	assign n_126 = ~n163;
	assign n_106 = ~n133;
	assign n_129 = ~n165;
	assign n407 = ( n_333 & n_139 );
	assign n223 = ( n_174 & n_175 );
	assign n_387 = ~n467;
	assign n489 = ( n_402 & n488 );
	assign n591 = ( n_491 & n_492 );
	assign n_63 = ~n80;
	assign n_80 = ~n101;
	assign n_608 = ~n137;
	assign n_288 = ~n358;
	assign n_427 = ~n517;
	assign n_211 = ~n264;
	assign n_241 = ~n303;
	assign n365 = ( n_118 & n_292 );
	assign n_363 = ~n440;
	assign n455 = ( n449 & n_375 );
	assign n495 = ( n_405 & n_406 );
	assign n_486 = ~n584;
	assign n_508 = ~n611;
	assign n123 = ( n_96 & n_97 );
	assign n182 = ( n_139 & n_140 );
	assign n_339 = ~n411;
	assign n664 = ( n_553 & n_554 );
	assign n_74 = ~n93;
	assign n_103 = ~n129;
	assign n_116 = ~n152;
	assign n_431 = ~n521;
	assign n_575 = ~n689;
	assign n_186 = ~n237;
	assign n_434 = ~n524;
	assign n_262 = ~n327;
	assign n_412 = ~n500;
	assign n_20 = ~n32;
	assign n468 = ( n_386 & n_387 );
	assign n600 = ( n_498 & n_499 );
	assign n_609 = ~n250;
	assign n638 = ( n_528 & n637 );
	assign n_70 = ~n88;
	assign n_305 = ~n194;
	assign n_494 = ~n305;
	assign n_238 = ~n300;
	assign n316 = ( n_249 & n_250 );
	assign n_269 = ~n334;
	assign n_373 = ~n450;
	assign n_470 = ~n566;
	assign n_521 = ~n628;
	assign n389 = ( n_316 & n388 );
	assign n_43 = ~n54;
	assign n_449 = ~n540;
	assign n_189 = ~n239;
	assign n_332 = ~n405;
	assign n_280 = ~n344;
	assign n_90 = ~n114;
	assign n_120 = ~n157;
	assign n_278 = ~n340;
	assign n_348 = ~n420;
	assign n_385 = ~n466;
	assign n_452 = ~n544;
	assign n_497 = ~n597;
	assign n_513 = ~n618;
	assign n_67 = ~n86;
	assign n_50 = ~n66;
	assign n_113 = ~n148;
	assign n_382 = ~n463;
	assign n_275 = ~n338;
	assign n_517 = ~n623;
	assign n_398 = ~n483;
	assign n_393 = ~n477;
	assign n_243 = ~n306;
	assign n_150 = ~n190;
	assign n_164 = ~n208;
	assign n_224 = ~n280;
	assign n_304 = ~n375;
	assign n_509 = ~n615;
	assign n_552 = ~n661;
	assign n_235 = ~n297;
	assign n_380 = ~n460;
	assign n_198 = ~n248;
	assign n_35 = ~n47;
	assign n_40 = ~n49;
	assign n_144 = ~n184;
	assign n_340 = ~n412;
	assign n_418 = ~n508;
	assign n_448 = ~n538;
	assign n_482 = ~n580;
	assign n_572 = ~n686;
	assign n_549 = ~n658;
	assign n_354 = ~n427;
	assign n33 = ( n_19 & n_20 );
	assign n_55 = ~n68;
	assign n_192 = ~n241;
	assign n_320 = ~n393;
	assign n_425 = ~n513;
	assign n_444 = ~n534;
	assign n_479 = ~n576;
	assign n_566 = ~n679;
	assign n_541 = ~n651;
	assign n_358 = ~n432;
	assign n_132 = ~n168;
	assign n_291 = ~n361;
	assign n_334 = ~n407;
	assign n_176 = ~n223;
	assign n_403 = ~n489;
	assign n_493 = ~n591;
	assign n_293 = ~n365;
	assign n_376 = ~n455;
	assign n_407 = ~n495;
	assign n_100 = ~n123;
	assign n_141 = ~n182;
	assign n_555 = ~n664;
	assign n_388 = ~n468_key;
	assign n_500 = ~n600_key;
	assign n_529 = ~n638_key;
	assign n_251 = ~n316_key;
	assign n_317 = ~n389_key;
	assign n_23 = ~n33_key;
	assign n33_key = ~( n33 ^ key_0 );
	assign n389_key = ~( n389 ^ key_1 );
	assign n316_key = ~( n316 ^ key_2 );
	assign n638_key = ~( n638 ^ key_3 );
	assign n600_key = ~( n600 ^ key_4 );
	assign n468_key = ~( n468 ^ key_5 );
	assign n317_key = ~( n317 ^ key_6 );
	assign n265_key = ~( n265 ^ key_7 );
	assign n275_key = ~( n275 ^ key_8 );
	assign n304_key = ~( n304 ^ key_9 );
	assign n345_key = ~( n345 ^ key_10 );
	assign n272_key = ~( n272 ^ key_11 );
	assign n307_key = ~( n307 ^ key_12 );
	assign n321_key = ~( n321 ^ key_13 );
	assign n262_key = ~( n262 ^ key_14 );
	assign n281_key = ~( n281 ^ key_15 );
	assign n328_key = ~( n328 ^ key_16 );
	assign n260_key = ~( n260 ^ key_17 );
	assign n274_key = ~( n274 ^ key_18 );
	assign n301_key = ~( n301 ^ key_19 );
	assign n311_key = ~( n311 ^ key_20 );
	assign n276_key = ~( n276 ^ key_21 );
	assign n323_key = ~( n323 ^ key_22 );
	assign n263_key = ~( n263 ^ key_23 );
	assign n314_key = ~( n314 ^ key_24 );
	assign n324_key = ~( n324 ^ key_25 );
	assign n331_key = ~( n331 ^ key_26 );
	assign n298_key = ~( n298 ^ key_27 );
	assign n346_key = ~( n346 ^ key_28 );
	assign n343_key = ~( n343 ^ key_29 );
	assign n337_key = ~( n337 ^ key_30 );
	assign n271_key = ~( n271 ^ key_31 );
	assign n279_key = ~( n279 ^ key_32 );
	assign n296_key = ~( n296 ^ key_33 );
	assign n284_key = ~( n284 ^ key_34 );
	assign n278_key = ~( n278 ^ key_35 );
	assign n312_key = ~( n312 ^ key_36 );
	assign n335_key = ~( n335 ^ key_37 );
	assign n302_key = ~( n302 ^ key_38 );
	assign n309_key = ~( n309 ^ key_39 );
	assign n289_key = ~( n289 ^ key_40 );
	assign n339_key = ~( n339 ^ key_41 );
	assign n350_key = ~( n350 ^ key_42 );
	assign n292_key = ~( n292 ^ key_43 );
	assign n258_key = ~( n258 ^ key_44 );
	assign n319_key = ~( n319 ^ key_45 );
	assign n341_key = ~( n341 ^ key_46 );
	assign n315_key = ~( n315 ^ key_47 );
	assign n270_key = ~( n270 ^ key_48 );
	assign n277_key = ~( n277 ^ key_49 );
	assign n318_key = ~( n318 ^ key_50 );
	assign n268_key = ~( n268 ^ key_51 );
	assign n330_key = ~( n330 ^ key_52 );
	assign n256_key = ~( n256 ^ key_53 );
	assign n269_key = ~( n269 ^ key_54 );
	assign n308_key = ~( n308 ^ key_55 );
	assign n347_key = ~( n347 ^ key_56 );
	assign n313_key = ~( n313 ^ key_57 );
	assign n273_key = ~( n273 ^ key_58 );
	assign n322_key = ~( n322 ^ key_59 );
	assign n326_key = ~( n326 ^ key_60 );
	assign n333_key = ~( n333 ^ key_61 );
	assign n288_key = ~( n288 ^ key_62 );
endmodule
