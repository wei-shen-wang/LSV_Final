module c3540(N1, N107, N116, N124, N125, N128, N13, N132, N137, N143, N150, N159, N169, N179, N190, N20, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N33, N330, N343, N349, N350, N41, N45, N50, N58, N68, N77, N87, N97, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361);
	input N1, N107, N116, N124, N125, N128, N13, N132, N137, N143, N150, N159, N169, N179, N190, N20, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N33, N330, N343, N349, N350, N41, N45, N50, N58, N68, N77, N87, N97;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20;
	output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361;
	wire N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350, N1562, N2482, AND3_113_inw1, AND3_208_inw1, N913, N1331, NAND3_59_inw1, NAND3_240_inw1, NAND3_271_inw1, NAND4_241_inw1, N769, N1197, N1219, N1409, N793, AND3_148_inw1, NAND3_117_inw1, N786, N890, N892, N1581, N1586, N1589, N1592, N1597, N1600, N2486, N2487, N1325, NAND3_240_invw, NAND4_241_inw2, N794, N1117, N829, N2022, N2024, N2026, N2028, N2030, N2032, N2034, N2036, N1738, N1818, NAND3_59_invw, N820, N896, n_88, n_101, n_114, n_127, n_140, n_153, n_177, N832, N835, N1322, N3387, N3389, AND3_111_inw1, NAND3_117_invw, N839, N1520, N1792, N3216, N3225, N3234, N3243, N3252, N3261, N3270, AND3_371_inw1, N2348, N1251, N2133, N1870, N665, N1787, N1794, N3224, N3233, N3242, N3251, N3260, N3269, AND3_372_inw1, AND4_401_inw2, N1252, N1960, N1875, N679, N1729, N1789, N1796, N3232, N3241, N3250, N3259, N3268, AND3_373_inw1, N1253, N1267, N1727, N2134, N1880, N686, N1791, N1798, N3240, N3249, N3258, N3267, AND3_374_inw1, AND3_468_inw1, N1254, N2135, N1885, N702, N1714, N1793, N1800, N3248, N3257, N3266, N3275, AND3_375_inw1, N1255, N2136, N1890, N724, N1795, N1802, N3256, N3265, N3276, N3283, N3290, AND3_376_inw1, N1256, N1961, N2137, N1895, N736, N1797, N3264, N3277, N3284, N3291, N3298, N3305, AND3_377_inw1, N1257, N1730, N2138, N1900, N749, N1799, N2349, N3278, N3285, N3292, N3299, N3306, N3313, N3320, AND3_378_inw1, N1258, N2139, N1905, N763, N3207, N3214, N3215, N3213, N3222, N3223, N3212, N3221, N3230, N3231, N3211, N3220, N3229, N3238, N3239, N3210, N3219, N3228, N3237, N3246, N3247, N1788, N3209, N3218, N3227, N3236, N3245, N3254, N3255, N1790, N3208, N3217, N3226, N3235, N3244, N3253, N3262, N3263, AND3_931_inw1, AND3_937_inw1, AND3_941_inw1, AND3_945_inw1, AND3_951_inw1, AND3_955_inw1, AND3_1023_inw1, AND3_1034_inw1, N1179, AND3_932_inw1, AND3_938_inw1, AND3_942_inw1, AND3_946_inw1, AND3_952_inw1, AND3_956_inw1, AND3_1024_inw1, AND3_1035_inw1, n_73, g7_inw2, AND3_933_inw1, AND3_939_inw1, AND3_943_inw1, AND3_947_inw1, AND3_953_inw1, AND3_957_inw1, AND3_1025_inw1, AND3_1036_inw1, N1358, N1803, AND3_934_inw1, AND3_940_inw1, AND3_944_inw1, AND3_948_inw1, AND3_954_inw1, AND3_958_inw1, AND3_1026_inw1, AND3_1037_inw1, N889, N1909, N5215, AND3_323_inw1, N920, N1643, N1644, N2023, N1645, N2025, AND3_481_inw1, N1510, N1259, N1646, N2027, AND3_484_inw1, N1509, N1260, N1647, N2029, AND3_487_inw1, N1512, N1261, N1648, N2031, AND3_490_inw1, N1511, N1262, N1067, N1649, N2033, AND3_493_inw1, N1692, N1467, N1650, N2035, AND3_496_inw1, N1691, N1468, N768, N2037, AND3_499_inw1, N1694, N1469, AND3_502_inw1, N1693, N1470, AND3_482_inw1, AND3_494_inw1, AND3_497_inw1, N1801, N3271, N3286, N3293, N3300, N3307, N3314, N3321, N3328, N3279, N3294, N3301, N3308, N3315, N3322, N3329, N3287, N3302, N3309, N3316, N3323, N3330, N3295, N3310, N3317, N3324, N3331, N3303, N3318, N3325, N3332, N3311, N3326, N3333, N3319, N3334, N3327, N4186, N4242, N4387, N4493, N4549, N4772, AND3_1289_inw1, AND3_1356_inw1, AND3_1381_inw1, N4515, N1460, g44_inw1, g93_inw1, N1913, N1464, N2307, N2730, N2121, N2761, N1667, N1202, N2184, N1770, NAND3_271_invw, NAND4_241_invw, N1306, N4498, N1869, N1196, N1452, N1833, NAND3_272_inw1, N1809, N891, N1806, N1366, OR3_345_inw1, OR3_346_inw1, OR3_347_inw1, OR3_348_inw1, OR3_349_inw1, OR3_350_inw1, OR3_602_inw1, OR3_603_inw1, N1983, N1747, N1328, N1756, N1580, N1579, N1426, OR3_440_inw1, OR3_441_inw1, OR3_442_inw1, OR3_443_inw1, OR3_444_inw1, OR3_445_inw1, OR3_446_inw1, OR3_447_inw1, N2144, N2143, N2211, n_164, N914, N1850, N1815, NAND3_272_invw, n_83, n_96, n_109, n_122, n_135, n_148, n_172, N1401, g23_inw2, g39_inw2, g56_inw2, g72_inw2, g88_inw2, g105_inw2, g135_inw2, N1315, N2436, N1893, N3534, N3536, N1337, N1966, N2350, N2376, N2758, N1987, g94_inw1, g124_invw, n_94, n_107, n_134, n_121, n_79, N2068, N2478, AND4_170_inw1, N2325, NOR3_553_inw1, N2398, N2898, AND3_86_inw1, N1940, N1988, g115_inw1, g124_inw1, g28_invw, n_133, n_82, N2073, N2148, N2146, NOR3_936_inw1, N2899, N1263, N1989, g28_inw1, g100_inw1, g45_invw, g115_invw, n_120, N2078, AND4_170_inw2, AND4_401_inw1, N2328, NOR3_557_inw1, N2900, N1250, N2769, g45_inw1, g130_inw1, g77_invw, g100_invw, n_162, n_81, N2083, NOR3_560_inw1, N2901, N1505, N1947, N1990, g34_inw1, g77_inw1, g61_invw, g130_invw, n_151, N2088, AND4_171_inw1, N2331, NOR3_563_inw1, N2347, AND3_120_inw1, N1991, g51_inw1, g61_inw1, g12_invw, g34_invw, n_163, n_175, N2093, N2147, NOR3_950_inw1, N2351, N1264, g12_inw1, g83_inw1, n_152, n_99, g51_invw, N2098, AND4_171_inw2, N2334, NOR3_567_inw1, N2355, N1340, N2483, n_176, n_112, g83_invw, g67_inw1, N2103, NOR3_570_inw1, N1722, N2353, g110_inw1, n_160, n_159, n_144, n_147, n_168, n_158, n_171, n_92, n_146, n_95, n_105, N1986, g110_invw, n_170, n_108, n_131, N2768, g94_invw, n_118, N3407, N3423, N3431, N3439, N3455, N3463, N3645, N3664, N3410, N3426, N3434, N3442, N3458, N3466, N3648, N3667, n_74, N3383, N3413, N3429, N3437, N3445, N3461, N3469, N3651, N3670, N2185, N2188, N2197, N2200, N1353, N2206, N3414, N3430, N3438, N3446, N3462, N3470, N3652, N3671, N3172, N3682, N1912, N5231, N2238, N2239, N2417, N1715, N2240, N2420, N2241, N2425, N1718, N2242, N2430, N2243, N2435, N1933, N2244, N2438, N2245, N2443, N1936, N2448, N2418, N2439, n_149, n_100, n_138, g67_invw, g18_inw1, n_173, n_113, n_125, g18_invw, n_97, n_139, n_86, n_110, n_126, n_136, n_87, n_123, n_84, N4675, N4291, N4678, N4461, N4786, N4596, N4716, N4558, N4924, N4706, N4859, N4817, N4331, N4545, N4608, N4559, N4463, N4390, N4435, N3175, N3178, N3181, N3184, N3187, N3605, N3690, N1917, N5136, N1461, N5277, N5286, N2310, g8_inw2, g24_inw2, g40_inw2, g57_inw2, g73_inw2, g89_inw2, g106_inw2, g120_inw2, N4647, N4794, N4800, N4831, N4838, N4907, N4913, N4985, NOR3_1373_invw, N2419, N2422, N2427, N2432, N2437, N2440, N2445, N2450, N2043, N1673, N4921, N2764, N1821, N1761, N1873, NOR3_1373_inw1, N2633, N2230, N2194, N1812, N2203, NOR3_590_inw1, N2145, N2181, N2180, N2980, N3388, N3632, N3633, g119_inw2, N1824, g17_inw2, g33_inw2, g50_inw2, g66_inw2, g82_inw2, g99_inw2, g129_inw2, N3552, N3544, N3546, N3550, N3548, N3540, N3542, N1898, OR3_564_inw1, N2277, n_169, g33_inw1, g50_inw1, NOR3_553_invw, N1507, N2755, N2474, N3634, n_156, N2282, n_93, g82_inw1, NOR3_936_invw, N2374, n_143, N2287, n_106, n_161, g66_inw1, NOR3_557_invw, N2754, N2475, n_167, N1338, N3149, n_132, n_150, g119_inw1, g17_inw1, NOR3_560_invw, n_91, N1713, N2352, N2294, n_119, n_174, g105_inw1, NOR3_563_invw, N1508, N2757, N2476, N3206, N2299, n_80, n_98, g135_inw1, NOR3_950_invw, N2375, N3535, g39_inw1, n_111, NOR3_567_invw, N2756, N2477, N3712, N1343, NOR3_1517_inw1, g56_inw1, n_137, NOR3_570_invw, N1725, N3711, g114_inw2, g114_inw1, g99_inw1, N2270, n_157, g129_inw1, N3119, n_145, N3644, N3657, N3661, N3663, N3676, N3680, N3789, N3803, g5_inw2, N3471, OR3_997_inw1, OR3_998_inw1, OR3_999_inw1, OR3_1000_inw1, OR3_1001_inw1, OR3_1002_inw1, OR3_1074_inw1, OR3_1078_inw1, N2984, N2985, N2988, N2989, N2191, N2991, N4075, N3681, N4147, N3898, N3912, OR3_554_inw1, N2749, N2467, OR3_555_inw1, OR3_558_inw1, N2748, N2468, OR3_561_inw1, N2342, N2141, OR3_565_inw1, OR3_568_inw1, N2341, N2142, OR3_571_inw1, g88_inw1, n_124, g72_inw1, n_85, g23_inw1, N4711, N4636, N4717, N4641, N4818, N4748, N4757, N4677, N4946, N4897, N4895, N4860, N4468, N4589, N4644, N4650, N4788, N4602, N4708, N4507, N4076, N3685, N4077, N3687, N4078, N3689, N4079, N3693, N4080, N3694, N4094, N4151, N3906, N3809, N3812, N3815, N3818, N3916, N4056, N4091, N5193, N5114, N5128, OR4_1640_inw1, OR4_1640_inw2, N5278, N5285, N4350, N4341, N4344, N4347, N4475, N4472, N4335, N4338, NOR3_1430_inw1, NOR3_1479_inw1, NOR3_1533_inw1, NOR3_1549_inw1, NOR3_1539_inw1, NOR3_1551_inw1, NOR3_1531_inw1, NOR3_1556_inw1, N4588, N2656, N2659, N2670, N2681, N2692, N2697, N2710, N2723, NOR3_1517_invw, N2641, N2632, N2481, N4189, N4191, N4192, N4303, N2987, N2990, NOR3_590_invw, N2354, OR3_780_inw1, OR3_979_inw1, N2379, OR3_1063_inw1, OR3_1064_inw1, N3538, N2234, N3551, N3543, N3545, N3549, N3547, N3539, N3541, N3641, N3637, N3638, N3640, N3639, N3635, N3636, N2652, N1721, N2973, N3713, N3419, N2666, N2677, N2688, N2977, N3406, N3451, N3642, N2706, N3779, N2719, N3780, N3537, N3721, NAND4_1153_inw1, N3734, N3654, N3740, N3658, N3743, NAND4_1154_inw1, N3756, N3673, N3762, N3677, N3838, N3786, N3845, N3800, N3194, N3557, N3568, N3573, N3578, N3589, N3594, N3731, N3753, N2986, N4105, N4029, N4190, N4106, N3947, N2966, N2471, N4797, N4808, AND4_1488_inw1, N4775, N4916, AND4_1526_inw1, N4889, N4905, N4904, AND4_1526_inw2, N4968, AND4_1488_inw2, N4900, N4442, N4981, N4870, N4823, N4754, N4743, N4674, N4107, N4030, N4108, N4031, N4109, N4032, N4111, N4033, N4112, N4034, N4284, N4317, AND4_1316_inw1, N4194, N4110, N4446, N3920, N4325, NAND3_1318_invw, N4421, N4327, N4287, N4238, N4393, NAND3_1286_invw, N4013, N3948, N4283, N4322, N4528, NAND3_1284_invw, NAND4_1319_inw2, N4295, N5242, N5201, N5223, N5222, N5298, NOR3_1430_invw, NOR3_1479_invw, NOR3_1531_invw, NOR3_1533_invw, NOR3_1539_invw, NOR3_1549_invw, NOR3_1556_invw, NOR3_1551_invw, N4667, N3115, N3125, N3131, N3138, N3145, N3155, g5_inw1, N3161, N3168, N4965, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N4954, N4957, N4973, N5010, N5013, N5030, n_155, n_166, n_90, n_142, N3195, OR3_1012_inw1, N4193, N4195, N4196, N4304, N2648, N3834, N3628, n_154, N3415, N2662, N2673, N2684, N3775, N3776, n_104, N3447, n_130, N2702, n_117, N2715, n_78, AND4_1130_inw1, N3894, NAND3_1131_inw1, NAND4_1132_inw2, N4042, NAND4_1153_invw, AND4_1130_inw2, N4043, NAND3_1131_invw, N4046, NAND4_1132_inw1, AND4_1133_inw1, N3895, NAND3_1134_inw1, NAND4_1135_inw2, N4049, NAND4_1154_invw, AND4_1133_inw2, N4050, NAND3_1134_invw, N4051, NAND4_1135_inw1, N4113, N4122, N4705, N4146, N4572, NAND3_1318_inw1, NAND4_1319_inw1, N4252, NAND4_1339_inw1, N3706, N3196, N3705, N3627, N4930, N4872, N4901, N4829, N4950, N4951, N4982, N4928, N4953, N4926, N5007, N4868, N4969, N4902, AND4_1316_inw2, N4552, NAND3_1284_inw1, N4148, g93_inw2, N4487, N4149, N4555, N4150, N4319, N4329, NAND3_1286_inw1, N4152, g44_inw2, N4153, N4668, N4506, N4443, N4573, N4256, NAND3_1310_inw1, N4447, N4509, N4508, NAND3_1312_inw1, N4530, N4496, N4458, N4328, N4310, N4576, N4326, NAND4_1319_invw, N5254, N5340, N5344, N4730, N4880, N4991, N4999, N5021, N5055, N5085, N5061, n_75, g7_inw1, N5002, n_141, n_165, n_89, n_102, n_128, n_115, n_76, g106_inw1, g120_inw1, g24_inw1, g89_inw1, n_103, n_116, n_77, n_129, N3987, N3926, NAND4_1132_invw, N3992, N3930, N3932, NAND4_1135_invw, N3996, N3935, N4740, N4670, N4619, N4527, NAND4_1339_invw, N3773, N4906, N4983, N4970, N4593, N4599, N4511, N4704, N4629, N4630, N4623, NAND3_1310_invw, NAND4_1339_inw2, NAND3_1312_invw, N4640, N4733, N4562, N4635, N4448, AND3_1630_inw1, AND3_1631_inw1, N5266, N5360, N5350, AND4_1552_inw1, N5094, N4815, AND4_1573_inw1, N5196, N4944, AND4_1552_inw2, N5110, N5045, N5108, N5047, N5125, N5078, AND3_1574_inw1, AND4_1573_inw2, N5183, N5102, N5212, N5120, N5220, N5121, g40_inw1, g73_inw1, g57_inw1, g8_inw1, N4028, N4073, N3931, N4074, NAND4_1153_inw2, N3936, NAND4_1154_inw2, N4896, N4673, N4503, N3833, N4931, N4984, N4747, N4753, N4676, N4416, N4427, N4769, N4688, AND3_1635_inw1, AND3_1636_inw1, N5066, N5122, N5133, N5236, N5145, N5228, N4104, N4669, N4526, N4510, N4816, N5166, N5245, N5217, N5284, N5250, N5232, N5233, N5295, N5253, N4145, N5192, N5258, N5309, N5354, N5279, N5348, N5352, N5358, N5361;
	wire N5358_key, N5348_key, N5354_key, N5309_key, N5258_key, N5295_key, N5232_key, N5183_key, N5212_key, N5228_key, N5284_key, N5094_key, N5196_key, N5110_key, N5108_key, N5125_key, N5220_key, N5122_key, N5236_key, N5145_key, N5245_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20;
	assign N1562 = ( N1 & N1337 );
	assign N2482 = ( N1761 & N1 );
	assign AND3_113_inw1 = ~( N1 & N786 );
	assign AND3_208_inw1 = ~( N1 & N13 );
	assign N913 = ~( N1 & N13 );
	assign N1331 = ~( N1 & N786 );
	assign NAND3_59_inw1 = ~( N1 & N20 );
	assign NAND3_240_inw1 = ~( N1 & N13 );
	assign NAND3_271_inw1 = ~( N1 & N13 );
	assign NAND4_241_inw1 = ~( N1 & N786 );
	assign N769 = ~N1;
	assign N1197 = ( N794 | N1 );
	assign N1219 = ( N820 | N1 );
	assign N1409 = ( N1 | N1196 );
	assign N793 = ( N13 & N20 );
	assign AND3_148_inw1 = ~( N769 & N13 );
	assign NAND3_117_inw1 = ~( N13 & N794 );
	assign N786 = ~N13;
	assign N890 = ( N20 & N200 );
	assign N892 = ( N20 & N179 );
	assign N1581 = ( N1338 & N20 );
	assign N1586 = ( N686 & N20 );
	assign N1589 = ( N77 & N20 );
	assign N1592 = ( N1343 & N20 );
	assign N1597 = ( N749 & N20 );
	assign N1600 = ( N116 & N20 );
	assign N2486 = ( N2374 & N20 );
	assign N2487 = ( N2375 & N20 );
	assign N1325 = ~( AND3_113_inw1 | N20 );
	assign NAND3_240_invw = ~( NAND3_240_inw1 | N20 );
	assign NAND4_241_inw2 = ~( N20 & N832 );
	assign N794 = ~N20;
	assign N1117 = ( N820 | N20 );
	assign N829 = ( N33 & N41 );
	assign N2022 = ( N77 & N33 );
	assign N2024 = ( N87 & N33 );
	assign N2026 = ( N97 & N33 );
	assign N2028 = ( N107 & N33 );
	assign N2030 = ( N116 & N33 );
	assign N2032 = ( N283 & N33 );
	assign N2034 = ( N294 & N33 );
	assign N2036 = ( N303 & N33 );
	assign N1738 = ~( N1325 & N33 );
	assign N1818 = ~( N33 & N832 );
	assign NAND3_59_invw = ~( NAND3_59_inw1 | N33 );
	assign N820 = ~N33;
	assign N896 = ( N349 | N33 );
	assign n_88 = ( n_84 & N33 );
	assign n_101 = ( n_97 & N33 );
	assign n_114 = ( n_110 & N33 );
	assign n_127 = ( n_123 & N33 );
	assign n_140 = ( n_136 & N33 );
	assign n_153 = ( n_149 & N33 );
	assign n_177 = ( n_173 & N33 );
	assign N832 = ~N41;
	assign N835 = ( N41 | N45 );
	assign N1322 = ( N769 & N45 );
	assign N3387 = ( N3196 & N45 );
	assign N3389 = ( N2973 & N45 );
	assign AND3_111_inw1 = ~( N769 & N45 );
	assign NAND3_117_invw = ~( NAND3_117_inw1 | N45 );
	assign N839 = ~N45;
	assign N1520 = ( N50 & N1263 );
	assign N1792 = ( N50 & N1580 );
	assign N3216 = ( N50 & N2985 );
	assign N3225 = ( N50 & N2986 );
	assign N3234 = ( N50 & N2987 );
	assign N3243 = ( N50 & N2988 );
	assign N3252 = ( N50 & N2989 );
	assign N3261 = ( N50 & N2990 );
	assign N3270 = ( N50 & N2991 );
	assign AND3_371_inw1 = ~( N50 & N1197 );
	assign N2348 = ~( AND3_468_inw1 | N50 );
	assign N1251 = ~( N226 & N50 );
	assign N2133 = ~( N50 & N58 );
	assign N1870 = ~( N50 | N1409 );
	assign N665 = ~N50;
	assign N1787 = ( N58 & N1579 );
	assign N1794 = ( N58 & N1580 );
	assign N3224 = ( N58 & N2985 );
	assign N3233 = ( N58 & N2986 );
	assign N3242 = ( N58 & N2987 );
	assign N3251 = ( N58 & N2988 );
	assign N3260 = ( N58 & N2989 );
	assign N3269 = ( N58 & N2990 );
	assign AND3_372_inw1 = ~( N58 & N1197 );
	assign AND4_401_inw2 = ~( N665 & N58 );
	assign N1252 = ~( N232 & N58 );
	assign N1960 = ~( N58 & N686 );
	assign N1875 = ~( N58 | N1409 );
	assign N679 = ~N58;
	assign N1729 = ( N68 & N665 );
	assign N1789 = ( N68 & N1579 );
	assign N1796 = ( N68 & N1580 );
	assign N3232 = ( N68 & N2985 );
	assign N3241 = ( N68 & N2986 );
	assign N3250 = ( N68 & N2987 );
	assign N3259 = ( N68 & N2988 );
	assign N3268 = ( N68 & N2989 );
	assign AND3_373_inw1 = ~( N68 & N1197 );
	assign N1253 = ~( N238 & N68 );
	assign N1267 = ~( N68 & N77 );
	assign N1727 = ~( N68 & N679 );
	assign N2134 = ~( N702 & N68 );
	assign N1880 = ~( N68 | N1409 );
	assign N686 = ~N68;
	assign N1791 = ( N77 & N1579 );
	assign N1798 = ( N77 & N1580 );
	assign N3240 = ( N77 & N2985 );
	assign N3249 = ( N77 & N2986 );
	assign N3258 = ( N77 & N2987 );
	assign N3267 = ( N77 & N2988 );
	assign AND3_374_inw1 = ~( N77 & N1197 );
	assign AND3_468_inw1 = ~( N2146 & N77 );
	assign N1254 = ~( N244 & N77 );
	assign N2135 = ~( N686 & N77 );
	assign N1885 = ~( N77 | N1409 );
	assign N702 = ~N77;
	assign N1714 = ( N87 & N1264 );
	assign N1793 = ( N87 & N1579 );
	assign N1800 = ( N87 & N1580 );
	assign N3248 = ( N87 & N2985 );
	assign N3257 = ( N87 & N2986 );
	assign N3266 = ( N87 & N2987 );
	assign N3275 = ( N87 & N2988 );
	assign AND3_375_inw1 = ~( N87 & N1219 );
	assign N1255 = ~( N250 & N87 );
	assign N2136 = ~( N736 & N87 );
	assign N1890 = ~( N87 | N1409 );
	assign N724 = ~N87;
	assign N1795 = ( N97 & N1579 );
	assign N1802 = ( N97 & N1580 );
	assign N3256 = ( N97 & N2985 );
	assign N3265 = ( N97 & N2986 );
	assign N3276 = ( N97 & N2989 );
	assign N3283 = ( N97 & N2988 );
	assign N3290 = ( N97 & N2987 );
	assign AND3_376_inw1 = ~( N97 & N1219 );
	assign N1256 = ~( N257 & N97 );
	assign N1961 = ~( N97 & N749 );
	assign N2137 = ~( N724 & N97 );
	assign N1895 = ~( N97 | N1409 );
	assign N736 = ~N97;
	assign N1797 = ( N107 & N1579 );
	assign N3264 = ( N107 & N2985 );
	assign N3277 = ( N107 & N2990 );
	assign N3284 = ( N107 & N2989 );
	assign N3291 = ( N107 & N2988 );
	assign N3298 = ( N107 & N2987 );
	assign N3305 = ( N107 & N2986 );
	assign AND3_377_inw1 = ~( N107 & N1219 );
	assign N1257 = ~( N264 & N107 );
	assign N1730 = ~( N107 & N736 );
	assign N2138 = ~( N763 & N107 );
	assign N1900 = ~( N107 | N1409 );
	assign N749 = ~N107;
	assign N1799 = ( N116 & N1579 );
	assign N2349 = ( N116 & N2147 );
	assign N3278 = ( N116 & N2991 );
	assign N3285 = ( N116 & N2990 );
	assign N3292 = ( N116 & N2989 );
	assign N3299 = ( N116 & N2988 );
	assign N3306 = ( N116 & N2987 );
	assign N3313 = ( N116 & N2986 );
	assign N3320 = ( N116 & N2985 );
	assign AND3_378_inw1 = ~( N116 & N1219 );
	assign N1258 = ~( N270 & N116 );
	assign N2139 = ~( N749 & N116 );
	assign N1905 = ~( N116 | N1409 );
	assign N763 = ~N116;
	assign N3207 = ( N124 & N2984 );
	assign N3214 = ( N125 & N2991 );
	assign N3215 = ( N125 & N2984 );
	assign N3213 = ( N128 & N2990 );
	assign N3222 = ( N128 & N2991 );
	assign N3223 = ( N128 & N2984 );
	assign N3212 = ( N132 & N2989 );
	assign N3221 = ( N132 & N2990 );
	assign N3230 = ( N132 & N2991 );
	assign N3231 = ( N132 & N2984 );
	assign N3211 = ( N137 & N2988 );
	assign N3220 = ( N137 & N2989 );
	assign N3229 = ( N137 & N2990 );
	assign N3238 = ( N137 & N2991 );
	assign N3239 = ( N137 & N2984 );
	assign N3210 = ( N143 & N2987 );
	assign N3219 = ( N143 & N2988 );
	assign N3228 = ( N143 & N2989 );
	assign N3237 = ( N143 & N2990 );
	assign N3246 = ( N143 & N2991 );
	assign N3247 = ( N143 & N2984 );
	assign N1788 = ( N150 & N1580 );
	assign N3209 = ( N150 & N2986 );
	assign N3218 = ( N150 & N2987 );
	assign N3227 = ( N150 & N2988 );
	assign N3236 = ( N150 & N2989 );
	assign N3245 = ( N150 & N2990 );
	assign N3254 = ( N150 & N2991 );
	assign N3255 = ( N150 & N2984 );
	assign N1790 = ( N159 & N1580 );
	assign N3208 = ( N159 & N2985 );
	assign N3217 = ( N159 & N2986 );
	assign N3226 = ( N159 & N2987 );
	assign N3235 = ( N159 & N2988 );
	assign N3244 = ( N159 & N2989 );
	assign N3253 = ( N159 & N2990 );
	assign N3262 = ( N159 & N2991 );
	assign N3263 = ( N159 & N2984 );
	assign AND3_931_inw1 = ~( N169 & N2648 );
	assign AND3_937_inw1 = ~( N169 & N2662 );
	assign AND3_941_inw1 = ~( N169 & N2673 );
	assign AND3_945_inw1 = ~( N169 & N2684 );
	assign AND3_951_inw1 = ~( N169 & N2702 );
	assign AND3_955_inw1 = ~( N169 & N2715 );
	assign AND3_1023_inw1 = ~( N169 & N3415 );
	assign AND3_1034_inw1 = ~( N169 & N3447 );
	assign N1179 = ( N794 | N169 );
	assign AND3_932_inw1 = ~( N179 & N2648 );
	assign AND3_938_inw1 = ~( N179 & N2662 );
	assign AND3_942_inw1 = ~( N179 & N2673 );
	assign AND3_946_inw1 = ~( N179 & N2684 );
	assign AND3_952_inw1 = ~( N179 & N2702 );
	assign AND3_956_inw1 = ~( N179 & N2715 );
	assign AND3_1024_inw1 = ~( N179 & N3415 );
	assign AND3_1035_inw1 = ~( N179 & N3447 );
	assign n_73 = ~N179;
	assign g7_inw2 = ~( N179 & n_75 );
	assign AND3_933_inw1 = ~( N190 & N2652 );
	assign AND3_939_inw1 = ~( N190 & N2666 );
	assign AND3_943_inw1 = ~( N190 & N2677 );
	assign AND3_947_inw1 = ~( N190 & N2688 );
	assign AND3_953_inw1 = ~( N190 & N2706 );
	assign AND3_957_inw1 = ~( N190 & N2719 );
	assign AND3_1025_inw1 = ~( N190 & N3419 );
	assign AND3_1036_inw1 = ~( N190 & N3451 );
	assign N1358 = ~( N794 | N190 );
	assign N1803 = ( N200 & N892 );
	assign AND3_934_inw1 = ~( N200 & N2652 );
	assign AND3_940_inw1 = ~( N200 & N2666 );
	assign AND3_944_inw1 = ~( N200 & N2677 );
	assign AND3_948_inw1 = ~( N200 & N2688 );
	assign AND3_954_inw1 = ~( N200 & N2706 );
	assign AND3_958_inw1 = ~( N200 & N2719 );
	assign AND3_1026_inw1 = ~( N200 & N3419 );
	assign AND3_1037_inw1 = ~( N200 & N3451 );
	assign N889 = ~N200;
	assign N1909 = ( N1452 & N213 );
	assign N5215 = ( N213 & N5193 );
	assign AND3_323_inw1 = ~( N1452 & N213 );
	assign N920 = ~N213;
	assign N1643 = ( N222 & N1401 );
	assign N1644 = ( N223 & N1401 );
	assign N2023 = ( N223 & N1850 );
	assign N1645 = ( N226 & N1401 );
	assign N2025 = ( N226 & N1850 );
	assign AND3_481_inw1 = ~( N2043 & N226 );
	assign N1510 = ~( N226 & N1260 );
	assign N1259 = ~N226;
	assign N1646 = ( N232 & N1401 );
	assign N2027 = ( N232 & N1850 );
	assign AND3_484_inw1 = ~( N2043 & N232 );
	assign N1509 = ~( N232 & N1259 );
	assign N1260 = ~N232;
	assign N1647 = ( N238 & N1401 );
	assign N2029 = ( N238 & N1850 );
	assign AND3_487_inw1 = ~( N2043 & N238 );
	assign N1512 = ~( N238 & N1262 );
	assign N1261 = ~N238;
	assign N1648 = ( N244 & N1401 );
	assign N2031 = ( N244 & N1850 );
	assign AND3_490_inw1 = ~( N2043 & N244 );
	assign N1511 = ~( N244 & N1261 );
	assign N1262 = ~N244;
	assign N1067 = ( N250 & N768 );
	assign N1649 = ( N250 & N1401 );
	assign N2033 = ( N250 & N1850 );
	assign AND3_493_inw1 = ~( N2043 & N250 );
	assign N1692 = ~( N250 & N1468 );
	assign N1467 = ~N250;
	assign N1650 = ( N257 & N1401 );
	assign N2035 = ( N257 & N1850 );
	assign AND3_496_inw1 = ~( N2043 & N257 );
	assign N1691 = ~( N257 & N1467 );
	assign N1468 = ~N257;
	assign N768 = ( N257 | N264 );
	assign N2037 = ( N264 & N1850 );
	assign AND3_499_inw1 = ~( N2043 & N264 );
	assign N1694 = ~( N264 & N1470 );
	assign N1469 = ~N264;
	assign AND3_502_inw1 = ~( N2043 & N270 );
	assign N1693 = ~( N270 & N1469 );
	assign N1470 = ~N270;
	assign AND3_482_inw1 = ~( N2043 & N274 );
	assign AND3_494_inw1 = ~( N2043 & N274 );
	assign AND3_497_inw1 = ~( N2043 & N274 );
	assign N1801 = ( N283 & N1579 );
	assign N3271 = ( N283 & N2984 );
	assign N3286 = ( N283 & N2991 );
	assign N3293 = ( N283 & N2990 );
	assign N3300 = ( N283 & N2989 );
	assign N3307 = ( N283 & N2988 );
	assign N3314 = ( N283 & N2987 );
	assign N3321 = ( N283 & N2986 );
	assign N3328 = ( N283 & N2985 );
	assign N3279 = ( N294 & N2984 );
	assign N3294 = ( N294 & N2991 );
	assign N3301 = ( N294 & N2990 );
	assign N3308 = ( N294 & N2989 );
	assign N3315 = ( N294 & N2988 );
	assign N3322 = ( N294 & N2987 );
	assign N3329 = ( N294 & N2986 );
	assign N3287 = ( N303 & N2984 );
	assign N3302 = ( N303 & N2991 );
	assign N3309 = ( N303 & N2990 );
	assign N3316 = ( N303 & N2989 );
	assign N3323 = ( N303 & N2988 );
	assign N3330 = ( N303 & N2987 );
	assign N3295 = ( N311 & N2984 );
	assign N3310 = ( N311 & N2991 );
	assign N3317 = ( N311 & N2990 );
	assign N3324 = ( N311 & N2989 );
	assign N3331 = ( N311 & N2988 );
	assign N3303 = ( N317 & N2984 );
	assign N3318 = ( N317 & N2991 );
	assign N3325 = ( N317 & N2990 );
	assign N3332 = ( N317 & N2989 );
	assign N3311 = ( N322 & N2984 );
	assign N3326 = ( N322 & N2991 );
	assign N3333 = ( N322 & N2990 );
	assign N3319 = ( N326 & N2984 );
	assign N3334 = ( N326 & N2991 );
	assign N3327 = ( N329 & N2984 );
	assign N4186 = ( N330 & N4094 );
	assign N4242 = ( N330 & N4112 );
	assign N4387 = ( N330 & N4317 );
	assign N4493 = ( N330 & N4319 );
	assign N4549 = ( N330 & N4443 );
	assign N4772 = ( N330 & N4704 );
	assign AND3_1289_inw1 = ~( N330 & N4094 );
	assign AND3_1356_inw1 = ~( N330 & N4319 );
	assign AND3_1381_inw1 = ~( N330 & N4284 );
	assign N4515 = ~( N330 & N4153 );
	assign N1460 = ~N330;
	assign g44_inw1 = ~( N330 & N4112 );
	assign g93_inw1 = ~( N330 & N4094 );
	assign N1913 = ~( AND3_323_inw1 | N343 );
	assign N1464 = ~( N920 | N343 );
	assign N2307 = ( N1464 & N350 );
	assign N2730 = ( N1562 & N1761 );
	assign N2121 = ~N1562;
	assign N2761 = ( N1722 & N2482 );
	assign N1667 = ~( AND3_208_inw1 | N1426 );
	assign N1202 = ( N913 & N914 );
	assign N2184 = ( N1331 & N1756 );
	assign N1770 = ~N1331;
	assign NAND3_271_invw = ~( NAND3_271_inw1 | N1179 );
	assign NAND4_241_invw = ~( NAND4_241_inw1 | NAND4_241_inw2 );
	assign N1306 = ( N769 & N835 );
	assign N4498 = ( N4442 & N769 );
	assign N1869 = ( N1202 & N1409 );
	assign N1196 = ~N793;
	assign N1452 = ~( AND3_148_inw1 | N794 );
	assign N1833 = ~( N786 & N820 );
	assign NAND3_272_inw1 = ~( N786 & N794 );
	assign N1809 = ( N890 & N1366 );
	assign N891 = ~N890;
	assign N1806 = ( N889 & N892 );
	assign N1366 = ~N892;
	assign OR3_345_inw1 = ~( N1581 | N1787 );
	assign OR3_346_inw1 = ~( N1586 | N1791 );
	assign OR3_347_inw1 = ~( N1589 | N1793 );
	assign OR3_348_inw1 = ~( N1592 | N1795 );
	assign OR3_349_inw1 = ~( N1597 | N1799 );
	assign OR3_350_inw1 = ~( N1600 | N1801 );
	assign OR3_602_inw1 = ~( N2486 | N1789 );
	assign OR3_603_inw1 = ~( N2487 | N1797 );
	assign N1983 = ( N1067 & N1325 );
	assign N1747 = ~( N1325 & N820 );
	assign N1328 = ~N1325;
	assign N1756 = ~NAND3_240_invw;
	assign N1580 = ( N794 & N1117 );
	assign N1579 = ~N1117;
	assign N1426 = ~N829;
	assign OR3_440_inw1 = ~( N2022 | N1643 );
	assign OR3_441_inw1 = ~( N2024 | N1644 );
	assign OR3_442_inw1 = ~( N2026 | N1645 );
	assign OR3_443_inw1 = ~( N2028 | N1646 );
	assign OR3_444_inw1 = ~( N2030 | N1647 );
	assign OR3_445_inw1 = ~( N2032 | N1648 );
	assign OR3_446_inw1 = ~( N2034 | N1649 );
	assign OR3_447_inw1 = ~( N2036 | N1650 );
	assign N2144 = ( N1738 & N1747 );
	assign N2143 = ~N1738;
	assign N2211 = ( N1815 & N1818 );
	assign n_164 = ~( N3278 | N1818 );
	assign N914 = ~NAND3_59_invw;
	assign N1850 = ( N820 & N896 );
	assign N1815 = ~( N820 & N832 );
	assign NAND3_272_invw = ~( NAND3_272_inw1 | N820 );
	assign n_83 = ( n_79 & N820 );
	assign n_96 = ( n_92 & N820 );
	assign n_109 = ( n_105 & N820 );
	assign n_122 = ( n_118 & N820 );
	assign n_135 = ( n_131 & N820 );
	assign n_148 = ( n_144 & N820 );
	assign n_172 = ( n_168 & N820 );
	assign N1401 = ~N896;
	assign g23_inw2 = ~( n_87 & n_88 );
	assign g39_inw2 = ~( n_100 & n_101 );
	assign g56_inw2 = ~( n_113 & n_114 );
	assign g72_inw2 = ~( n_126 & n_127 );
	assign g88_inw2 = ~( n_139 & n_140 );
	assign g105_inw2 = ~( n_152 & n_153 );
	assign g135_inw2 = ~( n_176 & n_177 );
	assign N1315 = ~( AND3_111_inw1 | N832 );
	assign N2436 = ~( AND3_494_inw1 | N1322 );
	assign N1893 = ~N1322;
	assign N3534 = ~( N3387 | N2350 );
	assign N3536 = ~( N3389 | N1966 );
	assign N1337 = ~NAND3_117_invw;
	assign N1966 = ( N1520 & N839 );
	assign N2350 = ( N2148 & N839 );
	assign N2376 = ( N1520 & N2180 );
	assign N2758 = ( N1520 & N2481 );
	assign N1987 = ~( OR3_346_inw1 & N1792 );
	assign g94_inw1 = ~( N3215 | N3216 );
	assign g124_invw = ~( g124_inw1 & N3225 );
	assign n_94 = ~( N3234 | N3235 );
	assign n_107 = ~( N3242 | N3243 );
	assign n_134 = ~( N3252 | N3253 );
	assign n_121 = ~( N3260 | N3261 );
	assign n_79 = ~N3270;
	assign N2068 = ~( AND3_371_inw1 | N1869 );
	assign N2478 = ( N2348 | N1729 );
	assign AND4_170_inw1 = ~( N1251 & N1252 );
	assign N2325 = ~( N1940 & N2133 );
	assign NOR3_553_inw1 = ~( N2270 | N1870 );
	assign N2398 = ( N665 & N2211 );
	assign N2898 = ( N665 & N2633 );
	assign AND3_86_inw1 = ~( N665 & N679 );
	assign N1940 = ~( N679 & N665 );
	assign N1988 = ~( OR3_347_inw1 & N1794 );
	assign g115_inw1 = ~( N3271 | N3224 );
	assign g124_inw1 = ~( N3223 | N3224 );
	assign g28_invw = ~( g28_inw1 & N3233 );
	assign n_133 = ~( N3250 | N3251 );
	assign n_82 = ~( N3268 | N3269 );
	assign N2073 = ~( AND3_372_inw1 | N1869 );
	assign N2148 = ~( AND4_401_inw1 | AND4_401_inw2 );
	assign N2146 = ~( N1727 & N1960 );
	assign NOR3_936_inw1 = ~( N3119 | N1875 );
	assign N2899 = ( N679 & N2633 );
	assign N1263 = ~( N679 & N686 );
	assign N1989 = ~( OR3_348_inw1 & N1796 );
	assign g28_inw1 = ~( N3231 | N3232 );
	assign g100_inw1 = ~( N3279 | N3232 );
	assign g45_invw = ~( g45_inw1 & N3241 );
	assign g115_invw = ~( g115_inw1 & N3241 );
	assign n_120 = ~( N3258 | N3259 );
	assign N2078 = ~( AND3_373_inw1 | N1869 );
	assign AND4_170_inw2 = ~( N1253 & N1254 );
	assign AND4_401_inw1 = ~( N1722 & N1267 );
	assign N2328 = ~( N2134 & N2135 );
	assign NOR3_557_inw1 = ~( N2277 | N1880 );
	assign N2900 = ( N686 & N2633 );
	assign N1250 = ~( AND3_86_inw1 | N686 );
	assign N2769 = ~( OR3_603_inw1 & N1798 );
	assign g45_inw1 = ~( N3239 | N3240 );
	assign g130_inw1 = ~( N3287 | N3240 );
	assign g77_invw = ~( g77_inw1 & N3249 );
	assign g100_invw = ~( g100_inw1 & N3249 );
	assign n_162 = ~( N3258 | N3275 );
	assign n_81 = ~( N3266 | N3267 );
	assign N2083 = ~( AND3_374_inw1 | N1869 );
	assign NOR3_560_inw1 = ~( N2282 | N1885 );
	assign N2901 = ( N702 & N2633 );
	assign N1505 = ~( N702 & N1250 );
	assign N1947 = ~N1714;
	assign N1990 = ~( OR3_349_inw1 & N1800 );
	assign g34_inw1 = ~( N3295 | N3248 );
	assign g77_inw1 = ~( N3247 | N3248 );
	assign g61_invw = ~( g61_inw1 & N3257 );
	assign g130_invw = ~( g130_inw1 & N3257 );
	assign n_151 = ~( N3266 | N3283 );
	assign N2088 = ~( AND3_375_inw1 | N1869 );
	assign AND4_171_inw1 = ~( N1255 & N1256 );
	assign N2331 = ~( N2136 & N2137 );
	assign NOR3_563_inw1 = ~( N2287 | N1890 );
	assign N2347 = ( N724 & N2144 );
	assign AND3_120_inw1 = ~( N724 & N736 );
	assign N1991 = ~( OR3_350_inw1 & N1802 );
	assign g51_inw1 = ~( N3303 | N3256 );
	assign g61_inw1 = ~( N3255 | N3256 );
	assign g12_invw = ~( g12_inw1 & N3265 );
	assign g34_invw = ~( g34_inw1 & N3265 );
	assign n_163 = ~( N3276 | N3277 );
	assign n_175 = ~( N3290 | N3291 );
	assign N2093 = ~( AND3_376_inw1 | N1869 );
	assign N2147 = ~( N1730 & N1961 );
	assign NOR3_950_inw1 = ~( N3149 | N1895 );
	assign N2351 = ( N736 & N2144 );
	assign N1264 = ~( N736 & N749 );
	assign g12_inw1 = ~( N3263 | N3264 );
	assign g83_inw1 = ~( N3311 | N3264 );
	assign n_152 = ~( N3284 | N3285 );
	assign n_99 = ~( N3298 | N3299 );
	assign g51_invw = ~( g51_inw1 & N3305 );
	assign N2098 = ~( AND3_377_inw1 | N1869 );
	assign AND4_171_inw2 = ~( N1257 & N1258 );
	assign N2334 = ~( N2138 & N2139 );
	assign NOR3_567_inw1 = ~( N2294 | N1900 );
	assign N2355 = ( N749 & N2144 );
	assign N1340 = ~( AND3_120_inw1 | N749 );
	assign N2483 = ( N2349 & N2180 );
	assign n_176 = ~( N3292 | N3293 );
	assign n_112 = ~( N3306 | N3307 );
	assign g83_invw = ~( g83_inw1 & N3313 );
	assign g67_inw1 = ~( N3319 | N3320 );
	assign N2103 = ~( AND3_378_inw1 | N1869 );
	assign NOR3_570_inw1 = ~( N2299 | N1905 );
	assign N1722 = ( N763 & N1340 );
	assign N2353 = ( N763 & N2144 );
	assign g110_inw1 = ~( N3207 | N3208 );
	assign n_160 = ~( N3214 | N1815 );
	assign n_159 = ~( N3212 | N3213 );
	assign n_144 = ~N3222;
	assign n_147 = ~( N3220 | N3221 );
	assign n_168 = ~N3230;
	assign n_158 = ~( N3210 | N3211 );
	assign n_171 = ~( N3228 | N3229 );
	assign n_92 = ~N3238;
	assign n_146 = ~( N3218 | N3219 );
	assign n_95 = ~( N3236 | N3237 );
	assign n_105 = ~N3246;
	assign N1986 = ~( OR3_345_inw1 & N1788 );
	assign g110_invw = ~( g110_inw1 & N3209 );
	assign n_170 = ~( N3226 | N3227 );
	assign n_108 = ~( N3244 | N3245 );
	assign n_131 = ~N3254;
	assign N2768 = ~( OR3_602_inw1 & N1790 );
	assign g94_invw = ~( g94_inw1 & N3217 );
	assign n_118 = ~N3262;
	assign N3407 = ~( AND3_931_inw1 | N2656 );
	assign N3423 = ~( AND3_937_inw1 | N2670 );
	assign N3431 = ~( AND3_941_inw1 | N2681 );
	assign N3439 = ~( AND3_945_inw1 | N2692 );
	assign N3455 = ~( AND3_951_inw1 | N2710 );
	assign N3463 = ~( AND3_955_inw1 | N2723 );
	assign N3645 = ~( AND3_1023_inw1 | N2659 );
	assign N3664 = ~( AND3_1034_inw1 | N2697 );
	assign N3410 = ~( AND3_932_inw1 | N3115 );
	assign N3426 = ~( AND3_938_inw1 | N3131 );
	assign N3434 = ~( AND3_942_inw1 | N3138 );
	assign N3442 = ~( AND3_946_inw1 | N3145 );
	assign N3458 = ~( AND3_952_inw1 | N3161 );
	assign N3466 = ~( AND3_956_inw1 | N3168 );
	assign N3648 = ~( AND3_1024_inw1 | N3125 );
	assign N3667 = ~( AND3_1035_inw1 | N3155 );
	assign n_74 = ( n_73 & N2692 );
	assign N3383 = ~( g7_inw1 | g7_inw2 );
	assign N3413 = ~( AND3_933_inw1 | N3115 );
	assign N3429 = ~( AND3_939_inw1 | N3131 );
	assign N3437 = ~( AND3_943_inw1 | N3138 );
	assign N3445 = ~( AND3_947_inw1 | N3145 );
	assign N3461 = ~( AND3_953_inw1 | N3161 );
	assign N3469 = ~( AND3_957_inw1 | N3168 );
	assign N3651 = ~( AND3_1025_inw1 | N3125 );
	assign N3670 = ~( AND3_1036_inw1 | N3155 );
	assign N2185 = ~( N1358 & N1812 );
	assign N2188 = ~( N1358 & N1809 );
	assign N2197 = ~( N1358 & N1806 );
	assign N2200 = ~( N1358 & N1803 );
	assign N1353 = ~N1358;
	assign N2206 = ~( N1353 & N1803 );
	assign N3414 = ~( AND3_934_inw1 | N2656 );
	assign N3430 = ~( AND3_940_inw1 | N2670 );
	assign N3438 = ~( AND3_944_inw1 | N2681 );
	assign N3446 = ~( AND3_948_inw1 | N2692 );
	assign N3462 = ~( AND3_954_inw1 | N2710 );
	assign N3470 = ~( AND3_958_inw1 | N2723 );
	assign N3652 = ~( AND3_1026_inw1 | N2659 );
	assign N3671 = ~( AND3_1037_inw1 | N2697 );
	assign N3172 = ( N1909 & N2648 );
	assign N3682 = ( N1909 & N3415 );
	assign N1912 = ~N1909;
	assign N5231 = ~N5215;
	assign N2238 = ~( OR3_440_inw1 & N2023 );
	assign N2239 = ~( OR3_441_inw1 & N2025 );
	assign N2417 = ~( AND3_481_inw1 | N1873 );
	assign N1715 = ~( N1509 & N1510 );
	assign N2240 = ~( OR3_442_inw1 & N2027 );
	assign N2420 = ~( AND3_484_inw1 | N1873 );
	assign N2241 = ~( OR3_443_inw1 & N2029 );
	assign N2425 = ~( AND3_487_inw1 | N1873 );
	assign N1718 = ~( N1511 & N1512 );
	assign N2242 = ~( OR3_444_inw1 & N2031 );
	assign N2430 = ~( AND3_490_inw1 | N1873 );
	assign N2243 = ~( OR3_445_inw1 & N2033 );
	assign N2435 = ~( AND3_493_inw1 | N1893 );
	assign N1933 = ~( N1691 & N1692 );
	assign N2244 = ~( OR3_446_inw1 & N2035 );
	assign N2438 = ~( AND3_496_inw1 | N1898 );
	assign N2245 = ~( OR3_447_inw1 & N2037 );
	assign N2443 = ~( AND3_499_inw1 | N1898 );
	assign N1936 = ~( N1693 & N1694 );
	assign N2448 = ~( AND3_502_inw1 | N1898 );
	assign N2418 = ~( AND3_482_inw1 | N1306 );
	assign N2439 = ~( AND3_497_inw1 | N1315 );
	assign n_149 = ~N3286;
	assign n_100 = ~( N3300 | N3301 );
	assign n_138 = ~( N3314 | N3315 );
	assign g67_invw = ~( g67_inw1 & N3321 );
	assign g18_inw1 = ~( N3327 | N3328 );
	assign n_173 = ~N3294;
	assign n_113 = ~( N3308 | N3309 );
	assign n_125 = ~( N3322 | N3323 );
	assign g18_invw = ~( g18_inw1 & N3329 );
	assign n_97 = ~N3302;
	assign n_139 = ~( N3316 | N3317 );
	assign n_86 = ~( N3330 | N3331 );
	assign n_110 = ~N3310;
	assign n_126 = ~( N3324 | N3325 );
	assign n_136 = ~N3318;
	assign n_87 = ~( N3332 | N3333 );
	assign n_123 = ~N3326;
	assign n_84 = ~N3334;
	assign N4675 = ~( N4186 & N4635 );
	assign N4291 = ~N4186;
	assign N4678 = ~( N4242 & N4640 );
	assign N4461 = ~N4242;
	assign N4786 = ~( N4387 & N4747 );
	assign N4596 = ~N4387;
	assign N4716 = ~( N4493 & N4676 );
	assign N4558 = ~N4493;
	assign N4924 = ~( N4549 & N4896 );
	assign N4706 = ~N4549;
	assign N4859 = ~( N4772 & N4816 );
	assign N4817 = ~N4772;
	assign N4331 = ~( AND3_1289_inw1 | N4295 );
	assign N4545 = ~( AND3_1356_inw1 | N4496 );
	assign N4608 = ~( AND3_1381_inw1 | N4562 );
	assign N4559 = ~( N4463 & N4515 );
	assign N4463 = ~( N4112 & N1460 );
	assign N4390 = ~( g44_inw1 | g44_inw2 );
	assign N4435 = ~( g93_inw1 | g93_inw2 );
	assign N3175 = ( N1913 & N2662 );
	assign N3178 = ( N1913 & N2673 );
	assign N3181 = ( N1913 & N2684 );
	assign N3184 = ( N1913 & N2702 );
	assign N3187 = ( N1913 & N2715 );
	assign N3605 = ( N3471 & N1913 );
	assign N3690 = ( N1913 & N3447 );
	assign N1917 = ~N1913;
	assign N5136 = ~( AND3_1574_inw1 | N1464 );
	assign N1461 = ~N1464;
	assign N5277 = ~( AND3_1630_inw1 | N2307 );
	assign N5286 = ~( AND3_1636_inw1 | N2307 );
	assign N2310 = ~N2307;
	assign g8_inw2 = ~( n_78 & N2730 );
	assign g24_inw2 = ~( n_91 & N2730 );
	assign g40_inw2 = ~( n_104 & N2730 );
	assign g57_inw2 = ~( n_117 & N2730 );
	assign g73_inw2 = ~( n_130 & N2730 );
	assign g89_inw2 = ~( n_143 & N2730 );
	assign g106_inw2 = ~( n_156 & N2730 );
	assign g120_inw2 = ~( n_167 & N2730 );
	assign N4647 = ( N4559 & N2121 );
	assign N4794 = ( N4711 & N2121 );
	assign N4800 = ( N4717 & N2121 );
	assign N4831 = ( N4743 & N2121 );
	assign N4838 = ( N4757 & N2121 );
	assign N4907 = ( N4818 & N2121 );
	assign N4913 = ( N4823 & N2121 );
	assign N4985 = ( N4946 & N2121 );
	assign NOR3_1373_invw = ~( NOR3_1373_inw1 & N2761 );
	assign N2419 = ( N1667 & N2238 );
	assign N2422 = ( N1667 & N2239 );
	assign N2427 = ( N1667 & N2240 );
	assign N2432 = ( N1667 & N2241 );
	assign N2437 = ( N1667 & N2242 );
	assign N2440 = ( N1667 & N2243 );
	assign N2445 = ( N1667 & N2244 );
	assign N2450 = ( N1667 & N2245 );
	assign N2043 = ~N1667;
	assign N1673 = ~N1202;
	assign N4921 = ( N4895 & N2184 );
	assign N2764 = ( N2478 & N1770 );
	assign N1821 = ~NAND3_271_invw;
	assign N1761 = ~NAND4_241_invw;
	assign N1873 = ~N1306;
	assign NOR3_1373_inw1 = ~( N2758 | N4498 );
	assign N2633 = ( N1821 & N1833 );
	assign N2230 = ~N1833;
	assign N2194 = ~( N1353 & N1809 );
	assign N1812 = ( N891 & N1366 );
	assign N2203 = ~( N1353 & N1806 );
	assign NOR3_590_inw1 = ~( N2376 | N1983 );
	assign N2145 = ~N1747;
	assign N2181 = ( N1756 & N1328 );
	assign N2180 = ~N1756;
	assign N2980 = ( N2471 & N2143 );
	assign N3388 = ( N2977 & N2143 );
	assign N3632 = ( N3536 & N2143 );
	assign N3633 = ( N3534 & N2143 );
	assign g119_inw2 = ~( n_163 & n_164 );
	assign N1824 = ~NAND3_272_invw;
	assign g17_inw2 = ~( n_82 & n_83 );
	assign g33_inw2 = ~( n_95 & n_96 );
	assign g50_inw2 = ~( n_108 & n_109 );
	assign g66_inw2 = ~( n_121 & n_122 );
	assign g82_inw2 = ~( n_134 & n_135 );
	assign g99_inw2 = ~( n_147 & n_148 );
	assign g129_inw2 = ~( n_171 & n_172 );
	assign N3552 = ~( g23_inw1 | g23_inw2 );
	assign N3544 = ~( g39_inw1 | g39_inw2 );
	assign N3546 = ~( g56_inw1 | g56_inw2 );
	assign N3550 = ~( g72_inw1 | g72_inw2 );
	assign N3548 = ~( g88_inw1 | g88_inw2 );
	assign N3540 = ~( g105_inw1 | g105_inw2 );
	assign N3542 = ~( g135_inw1 | g135_inw2 );
	assign N1898 = ~N1315;
	assign OR3_564_inw1 = ~( N2435 | N2436 );
	assign N2277 = ( N1987 & N1673 );
	assign n_169 = ~g124_invw;
	assign g33_inw1 = ~( n_93 & n_94 );
	assign g50_inw1 = ~( n_106 & n_107 );
	assign NOR3_553_invw = ~( NOR3_553_inw1 & N2068 );
	assign N1507 = ~( AND4_170_inw1 | AND4_170_inw2 );
	assign N2755 = ~( N2325 & N2475 );
	assign N2474 = ~N2325;
	assign N3634 = ~( OR3_1012_inw1 & N2398 );
	assign n_156 = ~N2898;
	assign N2282 = ( N1988 & N1673 );
	assign n_93 = ~g28_invw;
	assign g82_inw1 = ~( n_132 & n_133 );
	assign NOR3_936_invw = ~( NOR3_936_inw1 & N2073 );
	assign N2374 = ~N2146;
	assign n_143 = ~N2899;
	assign N2287 = ( N1989 & N1673 );
	assign n_106 = ~g45_invw;
	assign n_161 = ~g115_invw;
	assign g66_inw1 = ~( n_119 & n_120 );
	assign NOR3_557_invw = ~( NOR3_557_inw1 & N2078 );
	assign N2754 = ~( N2328 & N2474 );
	assign N2475 = ~N2328;
	assign n_167 = ~N2900;
	assign N1338 = ~N1250;
	assign N3149 = ( N2769 & N1673 );
	assign n_132 = ~g77_invw;
	assign n_150 = ~g100_invw;
	assign g119_inw1 = ~( n_161 & n_162 );
	assign g17_inw1 = ~( n_80 & n_81 );
	assign NOR3_560_invw = ~( NOR3_560_inw1 & N2083 );
	assign n_91 = ~N2901;
	assign N1713 = ~N1505;
	assign N2352 = ( N1947 & N2145 );
	assign N2294 = ( N1990 & N1673 );
	assign n_119 = ~g61_invw;
	assign n_174 = ~g130_invw;
	assign g105_inw1 = ~( n_150 & n_151 );
	assign NOR3_563_invw = ~( NOR3_563_inw1 & N2088 );
	assign N1508 = ~( AND4_171_inw1 | AND4_171_inw2 );
	assign N2757 = ~( N2331 & N2477 );
	assign N2476 = ~N2331;
	assign N3206 = ~( OR3_780_inw1 & N2347 );
	assign N2299 = ( N1991 & N1673 );
	assign n_80 = ~g12_invw;
	assign n_98 = ~g34_invw;
	assign g135_inw1 = ~( n_174 & n_175 );
	assign NOR3_950_invw = ~( NOR3_950_inw1 & N2093 );
	assign N2375 = ~N2147;
	assign N3535 = ~( OR3_979_inw1 & N2351 );
	assign g39_inw1 = ~( n_98 & n_99 );
	assign n_111 = ~g51_invw;
	assign NOR3_567_invw = ~( NOR3_567_inw1 & N2098 );
	assign N2756 = ~( N2334 & N2476 );
	assign N2477 = ~N2334;
	assign N3712 = ~( OR3_1064_inw1 & N2355 );
	assign N1343 = ~N1340;
	assign NOR3_1517_inw1 = ~( N2764 | N2483 );
	assign g56_inw1 = ~( n_111 & n_112 );
	assign n_137 = ~g83_invw;
	assign NOR3_570_invw = ~( NOR3_570_inw1 & N2103 );
	assign N1725 = ~N1722;
	assign N3711 = ~( OR3_1063_inw1 & N2353 );
	assign g114_inw2 = ~( n_159 & n_160 );
	assign g114_inw1 = ~( n_157 & n_158 );
	assign g99_inw1 = ~( n_145 & n_146 );
	assign N2270 = ( N1986 & N1673 );
	assign n_157 = ~g110_invw;
	assign g129_inw1 = ~( n_169 & n_170 );
	assign N3119 = ( N2768 & N1673 );
	assign n_145 = ~g94_invw;
	assign N3644 = ~( N3407 | N3410 );
	assign N3657 = ~( N3423 | N3426 );
	assign N3661 = ~( N3431 | N3434 );
	assign N3663 = ~( N3439 | N3442 );
	assign N3676 = ~( N3455 | N3458 );
	assign N3680 = ~( N3463 | N3466 );
	assign N3789 = ~( N3645 | N3648 );
	assign N3803 = ~( N3664 | N3667 );
	assign g5_inw2 = ~( N2723 & n_74 );
	assign N3471 = ( N3194 | N3383 );
	assign OR3_997_inw1 = ~( N3413 | N3414 );
	assign OR3_998_inw1 = ~( N3429 | N3430 );
	assign OR3_999_inw1 = ~( N3437 | N3438 );
	assign OR3_1000_inw1 = ~( N3445 | N3446 );
	assign OR3_1001_inw1 = ~( N3461 | N3462 );
	assign OR3_1002_inw1 = ~( N3469 | N3470 );
	assign OR3_1074_inw1 = ~( N3651 | N3652 );
	assign OR3_1078_inw1 = ~( N3670 | N3671 );
	assign N2984 = ~N2185;
	assign N2985 = ~N2188;
	assign N2988 = ~N2197;
	assign N2989 = ~N2200;
	assign N2191 = ~( N1353 & N1812 );
	assign N2991 = ~N2206;
	assign N4075 = ~( N3172 & N4042 );
	assign N3681 = ~N3172;
	assign N4147 = ~( N3682 & N4113 );
	assign N3898 = ~N3682;
	assign N3912 = ( N3786 & N1912 );
	assign OR3_554_inw1 = ~( N2417 | N2418 );
	assign N2749 = ~( N1715 & N2468 );
	assign N2467 = ~N1715;
	assign OR3_555_inw1 = ~( N2420 | N2418 );
	assign OR3_558_inw1 = ~( N2425 | N2418 );
	assign N2748 = ~( N1718 & N2467 );
	assign N2468 = ~N1718;
	assign OR3_561_inw1 = ~( N2430 | N2418 );
	assign N2342 = ~( N1933 & N2142 );
	assign N2141 = ~N1933;
	assign OR3_565_inw1 = ~( N2438 | N2439 );
	assign OR3_568_inw1 = ~( N2443 | N2439 );
	assign N2341 = ~( N1936 & N2141 );
	assign N2142 = ~N1936;
	assign OR3_571_inw1 = ~( N2448 | N2439 );
	assign g88_inw1 = ~( n_137 & n_138 );
	assign n_124 = ~g67_invw;
	assign g72_inw1 = ~( n_124 & n_125 );
	assign n_85 = ~g18_invw;
	assign g23_inw1 = ~( n_85 & n_86 );
	assign N4711 = ~( N4675 & N4636 );
	assign N4636 = ~( N4576 & N4291 );
	assign N4717 = ~( N4678 & N4641 );
	assign N4641 = ~( N4458 & N4461 );
	assign N4818 = ~( N4786 & N4748 );
	assign N4748 = ~( N4593 & N4596 );
	assign N4757 = ~( N4716 & N4677 );
	assign N4677 = ~( N4623 & N4558 );
	assign N4946 = ~( N4924 & N4897 );
	assign N4897 = ~( N4740 & N4706 );
	assign N4895 = ~( N4859 & N4860 );
	assign N4860 = ~( N4769 & N4817 );
	assign N4468 = ~( N4331 | N4091 );
	assign N4589 = ( N4545 | N4287 );
	assign N4644 = ~( N4608 | N4310 );
	assign N4650 = ( N4559 & N2481 );
	assign N4788 = ~( N4390 & N4753 );
	assign N4602 = ~N4390;
	assign N4708 = ~( N4435 & N4673 );
	assign N4507 = ~N4435;
	assign N4076 = ~( N3175 & N4043 );
	assign N3685 = ~N3175;
	assign N4077 = ~( N3178 & N4046 );
	assign N3687 = ~N3178;
	assign N4078 = ~( N3181 & N4049 );
	assign N3689 = ~N3181;
	assign N4079 = ~( N3184 & N4050 );
	assign N3693 = ~N3184;
	assign N4080 = ~( N3187 & N4051 );
	assign N3694 = ~N3187;
	assign N4094 = ( N3605 | N4056 );
	assign N4151 = ~( N3690 & N4122 );
	assign N3906 = ~N3690;
	assign N3809 = ( N3654 & N1917 );
	assign N3812 = ( N3658 & N1917 );
	assign N3815 = ( N3673 & N1917 );
	assign N3818 = ( N3677 & N1917 );
	assign N3916 = ( N3800 & N1917 );
	assign N4056 = ( N3932 & N1917 );
	assign N4091 = ( N3996 & N1917 );
	assign N5193 = ~( N5136 | N5166 );
	assign N5114 = ( N5102 & N1461 );
	assign N5128 = ( N1461 & N5120 );
	assign OR4_1640_inw1 = ~( N5277 | N5285 );
	assign OR4_1640_inw2 = ~( N5278 | N5286 );
	assign N5278 = ~( AND3_1631_inw1 | N2310 );
	assign N5285 = ~( AND3_1635_inw1 | N2310 );
	assign N4350 = ~( g8_inw1 | g8_inw2 );
	assign N4341 = ~( g24_inw1 | g24_inw2 );
	assign N4344 = ~( g40_inw1 | g40_inw2 );
	assign N4347 = ~( g57_inw1 | g57_inw2 );
	assign N4475 = ~( g73_inw1 | g73_inw2 );
	assign N4472 = ~( g89_inw1 | g89_inw2 );
	assign N4335 = ~( g106_inw1 | g106_inw2 );
	assign N4338 = ~( g120_inw1 | g120_inw2 );
	assign NOR3_1430_inw1 = ~( N4647 | N4650 );
	assign NOR3_1479_inw1 = ~( N4794 | N4797 );
	assign NOR3_1533_inw1 = ~( N4800 | N4957 );
	assign NOR3_1549_inw1 = ~( N4831 | N5010 );
	assign NOR3_1539_inw1 = ~( N4838 | N4973 );
	assign NOR3_1551_inw1 = ~( N4907 | N5013 );
	assign NOR3_1531_inw1 = ~( N4913 | N4954 );
	assign NOR3_1556_inw1 = ~( N4985 | N5030 );
	assign N4588 = ~NOR3_1373_invw;
	assign N2656 = ~( OR3_554_inw1 & N2419 );
	assign N2659 = ~( OR3_555_inw1 & N2422 );
	assign N2670 = ~( OR3_558_inw1 & N2427 );
	assign N2681 = ~( OR3_561_inw1 & N2432 );
	assign N2692 = ~( OR3_564_inw1 & N2437 );
	assign N2697 = ~( OR3_565_inw1 & N2440 );
	assign N2710 = ~( OR3_568_inw1 & N2445 );
	assign N2723 = ~( OR3_571_inw1 & N2450 );
	assign NOR3_1517_invw = ~( NOR3_1517_inw1 & N4921 );
	assign N2641 = ( N1821 & N1824 );
	assign N2632 = ~N1821;
	assign N2481 = ~N1761;
	assign N4189 = ( N4146 & N2230 );
	assign N4191 = ( N4148 & N2230 );
	assign N4192 = ( N4149 & N2230 );
	assign N4303 = ( N4252 & N2230 );
	assign N2987 = ~N2194;
	assign N2990 = ~N2203;
	assign NOR3_590_invw = ~( NOR3_590_inw1 & N2379 );
	assign N2354 = ( N1725 & N2145 );
	assign OR3_780_inw1 = ~( N2980 | N2145 );
	assign OR3_979_inw1 = ~( N3388 | N2145 );
	assign N2379 = ( N1721 & N2181 );
	assign OR3_1063_inw1 = ~( N3632 | N2352 );
	assign OR3_1064_inw1 = ~( N3633 | N2354 );
	assign N3538 = ~( g119_inw1 | g119_inw2 );
	assign N2234 = ~N1824;
	assign N3551 = ~( g17_inw1 | g17_inw2 );
	assign N3543 = ~( g33_inw1 | g33_inw2 );
	assign N3545 = ~( g50_inw1 | g50_inw2 );
	assign N3549 = ~( g66_inw1 | g66_inw2 );
	assign N3547 = ~( g82_inw1 | g82_inw2 );
	assign N3539 = ~( g99_inw1 | g99_inw2 );
	assign N3541 = ~( g129_inw1 | g129_inw2 );
	assign N3641 = ( N3551 | N3552 );
	assign N3637 = ( N3543 | N3544 );
	assign N3638 = ( N3545 | N3546 );
	assign N3640 = ( N3549 | N3550 );
	assign N3639 = ( N3547 | N3548 );
	assign N3635 = ( N3539 | N3540 );
	assign N3636 = ( N3541 | N3542 );
	assign N2652 = ~NOR3_553_invw;
	assign N1721 = ~( N1507 & N1508 );
	assign N2973 = ~( N2754 & N2755 );
	assign N3713 = ( N3634 & N2632 );
	assign N3419 = ~NOR3_936_invw;
	assign N2666 = ~NOR3_557_invw;
	assign N2677 = ~NOR3_560_invw;
	assign N2688 = ~NOR3_563_invw;
	assign N2977 = ~( N2756 & N2757 );
	assign N3406 = ( N3206 & N2641 );
	assign N3451 = ~NOR3_950_invw;
	assign N3642 = ( N3535 & N2641 );
	assign N2706 = ~NOR3_567_invw;
	assign N3779 = ( N3712 & N2641 );
	assign N2719 = ~NOR3_570_invw;
	assign N3780 = ( N3711 & N2641 );
	assign N3537 = ~( g114_inw1 | g114_inw2 );
	assign N3721 = ( N3644 & N3557 );
	assign NAND4_1153_inw1 = ~( N3644 & N3894 );
	assign N3734 = ( N3657 & N3568 );
	assign N3654 = ~N3657;
	assign N3740 = ( N3661 & N3573 );
	assign N3658 = ~N3661;
	assign N3743 = ( N3663 & N3578 );
	assign NAND4_1154_inw1 = ~( N3663 & N3895 );
	assign N3756 = ( N3676 & N3589 );
	assign N3673 = ~N3676;
	assign N3762 = ( N3680 & N3594 );
	assign N3677 = ~N3680;
	assign N3838 = ( N3789 & N3731 );
	assign N3786 = ~N3789;
	assign N3845 = ( N3803 & N3753 );
	assign N3800 = ~N3803;
	assign N3194 = ~( g5_inw1 | g5_inw2 );
	assign N3557 = ~( OR3_997_inw1 & N2648 );
	assign N3568 = ~( OR3_998_inw1 & N2662 );
	assign N3573 = ~( OR3_999_inw1 & N2673 );
	assign N3578 = ~( OR3_1000_inw1 & N2684 );
	assign N3589 = ~( OR3_1001_inw1 & N2702 );
	assign N3594 = ~( OR3_1002_inw1 & N2715 );
	assign N3731 = ~( OR3_1074_inw1 & N3415 );
	assign N3753 = ~( OR3_1078_inw1 & N3447 );
	assign N2986 = ~N2191;
	assign N4105 = ~( N4075 & N4029 );
	assign N4029 = ~( N3721 & N3681 );
	assign N4190 = ~( N4147 & N4106 );
	assign N4106 = ~( N3838 & N3898 );
	assign N3947 = ~N3912;
	assign N2966 = ~( N2748 & N2749 );
	assign N2471 = ~( N2341 & N2342 );
	assign N4797 = ( N4711 & N2481 );
	assign N4808 = ( N4717 & N4468 );
	assign AND4_1488_inw1 = ~( N4717 & N4757 );
	assign N4775 = ~N4717;
	assign N4916 = ( N4818 & N4644 );
	assign AND4_1526_inw1 = ~( N4818 & N4743 );
	assign N4889 = ~N4818;
	assign N4905 = ~( N4757 & N4872 );
	assign N4904 = ~N4757;
	assign AND4_1526_inw2 = ~( N4946 & N4644 );
	assign N4968 = ~N4946;
	assign AND4_1488_inw2 = ~( N4823 & N4468 );
	assign N4900 = ~( N4868 | N4468 );
	assign N4442 = ~N4468;
	assign N4981 = ~( N4968 | N4644 );
	assign N4870 = ~N4644;
	assign N4823 = ~( N4788 & N4754 );
	assign N4754 = ~( N4599 & N4602 );
	assign N4743 = ~( N4708 & N4674 );
	assign N4674 = ~( N4619 & N4507 );
	assign N4107 = ~( N4076 & N4030 );
	assign N4030 = ~( N3734 & N3685 );
	assign N4108 = ~( N4077 & N4031 );
	assign N4031 = ~( N3740 & N3687 );
	assign N4109 = ~( N4078 & N4032 );
	assign N4032 = ~( N3743 & N3689 );
	assign N4111 = ~( N4079 & N4033 );
	assign N4033 = ~( N3756 & N3693 );
	assign N4112 = ~( N4080 & N4034 );
	assign N4034 = ~( N3762 & N3694 );
	assign N4284 = ( N4094 & N3926 );
	assign N4317 = ( N4094 & N4108 );
	assign AND4_1316_inw1 = ~( N4094 & N4190 );
	assign N4194 = ~( N4151 & N4110 );
	assign N4110 = ~( N3845 & N3906 );
	assign N4446 = ~( N4190 & N3809 );
	assign N3920 = ~N3809;
	assign N4325 = ~( N4107 & N3812 );
	assign NAND3_1318_invw = ~( NAND3_1318_inw1 | N3812 );
	assign N4421 = ( N3812 | N4322 );
	assign N4327 = ~( N4194 & N3815 );
	assign N4287 = ( N3815 | N4238 );
	assign N4238 = ( N4111 & N3818 );
	assign N4393 = ~( N3818 & N4152 );
	assign NAND3_1286_invw = ~( NAND3_1286_inw1 | N3818 );
	assign N4013 = ~N3818;
	assign N3948 = ~N3916;
	assign N4283 = ( N4091 & N3926 );
	assign N4322 = ( N4091 & N4108 );
	assign N4528 = ~( N4091 & N4149 );
	assign NAND3_1284_invw = ~( NAND3_1284_inw1 | N4091 );
	assign NAND4_1319_inw2 = ~( N4108 & N4091 );
	assign N4295 = ~N4091;
	assign N5242 = ~( N5114 & N5222 );
	assign N5201 = ~N5114;
	assign N5223 = ~( N5128 & N5201 );
	assign N5222 = ~N5128;
	assign N5298 = ~( OR4_1640_inw1 & OR4_1640_inw2 );
	assign NOR3_1430_invw = ~( NOR3_1430_inw1 & N4350 );
	assign NOR3_1479_invw = ~( NOR3_1479_inw1 & N4341 );
	assign NOR3_1531_invw = ~( NOR3_1531_inw1 & N4344 );
	assign NOR3_1533_invw = ~( NOR3_1533_inw1 & N4347 );
	assign NOR3_1539_invw = ~( NOR3_1539_inw1 & N4475 );
	assign NOR3_1549_invw = ~( NOR3_1549_inw1 & N4472 );
	assign NOR3_1556_invw = ~( NOR3_1556_inw1 & N4335 );
	assign NOR3_1551_invw = ~( NOR3_1551_inw1 & N4338 );
	assign N4667 = ~N4588;
	assign N3115 = ~N2656;
	assign N3125 = ~N2659;
	assign N3131 = ~N2670;
	assign N3138 = ~N2681;
	assign N3145 = ~N2692;
	assign N3155 = ~N2697;
	assign g5_inw1 = ~( N2697 & N2710 );
	assign N3161 = ~N2710;
	assign N3168 = ~N2723;
	assign N4965 = ~NOR3_1517_invw;
	assign N3714 = ( N3635 & N2632 );
	assign N3715 = ( N3636 & N2632 );
	assign N3716 = ( N3637 & N2632 );
	assign N3717 = ( N3638 & N2632 );
	assign N3718 = ( N3639 & N2632 );
	assign N3719 = ( N3640 & N2632 );
	assign N3720 = ( N3641 & N2632 );
	assign N4954 = ( N4926 & N2481 );
	assign N4957 = ( N4931 & N2481 );
	assign N4973 = ( N4953 & N2481 );
	assign N5010 = ( N4983 & N2481 );
	assign N5013 = ( N4984 & N2481 );
	assign N5030 = ( N5007 & N2481 );
	assign n_155 = ~N4189;
	assign n_166 = ~N4191;
	assign n_90 = ~N4192;
	assign n_142 = ~N4303;
	assign N3195 = ~NOR3_590_invw;
	assign OR3_1012_inw1 = ~( N3537 | N3538 );
	assign N4193 = ( N4150 & N2234 );
	assign N4195 = ( N4152 & N2234 );
	assign N4196 = ( N4153 & N2234 );
	assign N4304 = ( N4256 & N2234 );
	assign N2648 = ~N2652;
	assign N3834 = ~( N2973 & N3776 );
	assign N3628 = ~N2973;
	assign n_154 = ~N3713;
	assign N3415 = ~N3419;
	assign N2662 = ~N2666;
	assign N2673 = ~N2677;
	assign N2684 = ~N2688;
	assign N3775 = ~( N2977 & N3628 );
	assign N3776 = ~N2977;
	assign n_104 = ~N3406;
	assign N3447 = ~N3451;
	assign n_130 = ~N3642;
	assign N2702 = ~N2706;
	assign n_117 = ~N3779;
	assign N2715 = ~N2719;
	assign n_78 = ~N3780;
	assign AND4_1130_inw1 = ~( N3721 & N3838 );
	assign N3894 = ~( N3721 & N3786 );
	assign NAND3_1131_inw1 = ~( N3721 & N3838 );
	assign NAND4_1132_inw2 = ~( N3734 & N3721 );
	assign N4042 = ~N3721;
	assign NAND4_1153_invw = ~( NAND4_1153_inw1 | NAND4_1153_inw2 );
	assign AND4_1130_inw2 = ~( N3734 & N3740 );
	assign N4043 = ~N3734;
	assign NAND3_1131_invw = ~( NAND3_1131_inw1 | N3654 );
	assign N4046 = ~N3740;
	assign NAND4_1132_inw1 = ~( N3658 & N3838 );
	assign AND4_1133_inw1 = ~( N3743 & N3845 );
	assign N3895 = ~( N3743 & N3800 );
	assign NAND3_1134_inw1 = ~( N3743 & N3845 );
	assign NAND4_1135_inw2 = ~( N3756 & N3743 );
	assign N4049 = ~N3743;
	assign NAND4_1154_invw = ~( NAND4_1154_inw1 | NAND4_1154_inw2 );
	assign AND4_1133_inw2 = ~( N3756 & N3762 );
	assign N4050 = ~N3756;
	assign NAND3_1134_invw = ~( NAND3_1134_inw1 | N3673 );
	assign N4051 = ~N3762;
	assign NAND4_1135_inw1 = ~( N3677 & N3845 );
	assign N4113 = ~N3838;
	assign N4122 = ~N3845;
	assign N4705 = ~( N4105 & N4669 );
	assign N4146 = ~N4105;
	assign N4572 = ~( N4190 & N4526 );
	assign NAND3_1318_inw1 = ~( N4190 & N4107 );
	assign NAND4_1319_inw1 = ~( N4190 & N4107 );
	assign N4252 = ~N4190;
	assign NAND4_1339_inw1 = ~( N3947 & N4446 );
	assign N3706 = ~( N2966 & N3627 );
	assign N3196 = ~N2966;
	assign N3705 = ~( N2471 & N3196 );
	assign N3627 = ~N2471;
	assign N4930 = ~( N4808 & N4904 );
	assign N4872 = ~N4808;
	assign N4901 = ~( AND4_1488_inw1 | AND4_1488_inw2 );
	assign N4829 = ~( N4775 & N4442 );
	assign N4950 = ~( N4916 & N4902 );
	assign N4951 = ~N4916;
	assign N4982 = ~( AND4_1526_inw1 | AND4_1526_inw2 );
	assign N4928 = ~( N4889 & N4870 );
	assign N4953 = ~( N4930 & N4905 );
	assign N4926 = ( N4900 | N4901 );
	assign N5007 = ( N4981 | N4982 );
	assign N4868 = ~N4823;
	assign N4969 = ~( N4743 & N4951 );
	assign N4902 = ~N4743;
	assign AND4_1316_inw2 = ~( N4107 & N4108 );
	assign N4552 = ~( N4107 & N4508 );
	assign NAND3_1284_inw1 = ~( N4107 & N4108 );
	assign N4148 = ~N4107;
	assign g93_inw2 = ~( N4108 & N4107 );
	assign N4487 = ~( N4108 & N4295 );
	assign N4149 = ~N4108;
	assign N4555 = ~( N4109 & N4510 );
	assign N4150 = ~N4109;
	assign N4319 = ( N4112 & N4111 );
	assign N4329 = ~( N4111 & N4013 );
	assign NAND3_1286_inw1 = ~( N4194 & N4111 );
	assign N4152 = ~N4111;
	assign g44_inw2 = ~( N4111 & N4194 );
	assign N4153 = ~N4112;
	assign N4668 = ~( N4284 & N4630 );
	assign N4506 = ~N4284;
	assign N4443 = ~( AND4_1316_inw1 | AND4_1316_inw2 );
	assign N4573 = ~( N4194 & N4496 );
	assign N4256 = ~N4194;
	assign NAND3_1310_inw1 = ~( N3920 & N4325 );
	assign N4447 = ~NAND3_1318_invw;
	assign N4509 = ~( N4421 & N4148 );
	assign N4508 = ~N4421;
	assign NAND3_1312_inw1 = ~( N3948 & N4327 );
	assign N4530 = ~( N4287 & N4256 );
	assign N4496 = ~N4287;
	assign N4458 = ~( N4329 & N4393 );
	assign N4328 = ~NAND3_1286_invw;
	assign N4310 = ( N3992 | N4283 );
	assign N4576 = ~( N4487 & N4528 );
	assign N4326 = ~NAND3_1284_invw;
	assign NAND4_1319_invw = ~( NAND4_1319_inw1 | NAND4_1319_inw2 );
	assign N5254 = ~( N5242 & N5223 );
	assign N5340 = ~( N5298 & N5258_key );
	assign N5344 = ~N5298;
	assign N4730 = ~NOR3_1430_invw;
	assign N4880 = ~NOR3_1479_invw;
	assign N4991 = ~NOR3_1531_invw;
	assign N4999 = ~NOR3_1533_invw;
	assign N5021 = ~NOR3_1539_invw;
	assign N5055 = ~NOR3_1549_invw;
	assign N5085 = ~NOR3_1556_invw;
	assign N5061 = ~NOR3_1551_invw;
	assign n_75 = ( N3145 & N3155 );
	assign g7_inw1 = ~( N3161 & N3168 );
	assign N5002 = ~N4965;
	assign n_141 = ~N3714;
	assign n_165 = ~N3715;
	assign n_89 = ~N3716;
	assign n_102 = ~N3717;
	assign n_128 = ~N3718;
	assign n_115 = ~N3719;
	assign n_76 = ~N3720;
	assign g106_inw1 = ~( n_154 & n_155 );
	assign g120_inw1 = ~( n_165 & n_166 );
	assign g24_inw1 = ~( n_89 & n_90 );
	assign g89_inw1 = ~( n_141 & n_142 );
	assign n_103 = ~N4193;
	assign n_116 = ~N4195;
	assign n_77 = ~N4196;
	assign n_129 = ~N4304;
	assign N3987 = ~( N3775 & N3834 );
	assign N3926 = ~( AND4_1130_inw1 | AND4_1130_inw2 );
	assign NAND4_1132_invw = ~( NAND4_1132_inw1 | NAND4_1132_inw2 );
	assign N3992 = ~NAND4_1153_invw;
	assign N3930 = ~NAND3_1131_invw;
	assign N3932 = ~( AND4_1133_inw1 | AND4_1133_inw2 );
	assign NAND4_1135_invw = ~( NAND4_1135_inw1 | NAND4_1135_inw2 );
	assign N3996 = ~NAND4_1154_invw;
	assign N3935 = ~NAND3_1134_invw;
	assign N4740 = ~( N4705 & N4670 );
	assign N4670 = ~( N4503 & N4146 );
	assign N4619 = ~( N4572 & N4527 );
	assign N4527 = ~( N4416 & N4252 );
	assign NAND4_1339_invw = ~( NAND4_1339_inw1 | NAND4_1339_inw2 );
	assign N3773 = ~( N3705 & N3706 );
	assign N4906 = ~( N4872 & N4829 );
	assign N4983 = ~( N4950 & N4969 );
	assign N4970 = ~( N4951 & N4928 );
	assign N4593 = ~( N4552 & N4509 );
	assign N4599 = ~( N4555 & N4511 );
	assign N4511 = ~( N4427 & N4150 );
	assign N4704 = ~( N4629 & N4668 );
	assign N4629 = ~( N4443 & N4506 );
	assign N4630 = ~N4443;
	assign N4623 = ~( N4573 & N4530 );
	assign NAND3_1310_invw = ~( NAND3_1310_inw1 | N4326 );
	assign NAND4_1339_inw2 = ~( N4447 & N4448 );
	assign NAND3_1312_invw = ~( NAND3_1312_inw1 | N4328 );
	assign N4640 = ~N4458;
	assign N4733 = ~( N4310 & N4669 );
	assign N4562 = ~N4310;
	assign N4635 = ~N4576;
	assign N4448 = ~NAND4_1319_invw;
	assign AND3_1630_inw1 = ~( N5236_key & N5254 );
	assign AND3_1631_inw1 = ~( N5250 & N5254 );
	assign N5266 = ~N5254;
	assign N5360 = ~( N5350 & N5340 );
	assign N5350 = ~( N5279 & N5344 );
	assign AND4_1552_inw1 = ~( N4730 & N4999 );
	assign N5094 = ~( N5047 & N4730 );
	assign N4815 = ~N4730;
	assign AND4_1573_inw1 = ~( N4880 & N5061 );
	assign N5196 = ~( N5121 & N4880 );
	assign N4944 = ~N4880;
	assign AND4_1552_inw2 = ~( N5021 & N4991 );
	assign N5110 = ~( N5078 & N4991 );
	assign N5045 = ~N4991;
	assign N5108 = ~( N4815 & N4999 );
	assign N5047 = ~N4999;
	assign N5125 = ~( N5045 & N5021 );
	assign N5078 = ~N5021;
	assign AND3_1574_inw1 = ~( N5055 & N5085 );
	assign AND4_1573_inw2 = ~( N5055 & N5085 );
	assign N5183 = ~( N5120 & N5055 );
	assign N5102 = ~N5055;
	assign N5212 = ~( N5102 & N5085 );
	assign N5120 = ~N5085;
	assign N5220 = ~( N4944 & N5061 );
	assign N5121 = ~N5061;
	assign g40_inw1 = ~( n_102 & n_103 );
	assign g73_inw1 = ~( n_128 & n_129 );
	assign g57_inw1 = ~( n_115 & n_116 );
	assign g8_inw1 = ~( n_76 & n_77 );
	assign N4028 = ( N3932 & N3926 );
	assign N4073 = ~( N3926 & N3996 );
	assign N3931 = ~NAND4_1132_invw;
	assign N4074 = ~N3992;
	assign NAND4_1153_inw2 = ~( N3930 & N3931 );
	assign N3936 = ~NAND4_1135_invw;
	assign NAND4_1154_inw2 = ~( N3935 & N3936 );
	assign N4896 = ~N4740;
	assign N4673 = ~N4619;
	assign N4503 = ~NAND4_1339_invw;
	assign N3833 = ~N3773;
	assign N4931 = ~N4906;
	assign N4984 = ~N4970;
	assign N4747 = ~N4593;
	assign N4753 = ~N4599;
	assign N4676 = ~N4623;
	assign N4416 = ~NAND3_1310_invw;
	assign N4427 = ~NAND3_1312_invw;
	assign N4769 = ~( N4733 & N4688 );
	assign N4688 = ~( N4503 & N4562 );
	assign AND3_1635_inw1 = ~( N5236_key & N5266 );
	assign AND3_1636_inw1 = ~( N5250 & N5266 );
	assign N5066 = ~( AND4_1552_inw1 | AND4_1552_inw2 );
	assign N5122 = ~( N5094_key & N5108_key );
	assign N5133 = ~( AND4_1573_inw1 | AND4_1573_inw2 );
	assign N5236 = ~( N5196_key & N5220_key );
	assign N5145 = ~( N5125_key & N5110_key );
	assign N5228 = ~( N5183_key & N5212_key );
	assign N4104 = ( N4073 & N4074 );
	assign N4669 = ~N4503;
	assign N4526 = ~N4416;
	assign N4510 = ~N4427;
	assign N4816 = ~N4769;
	assign N5166 = ( N5066 & N5133 );
	assign N5245 = ~( N5122_key & N5233 );
	assign N5217 = ~N5122_key;
	assign N5284 = ~( N5236_key & N5253 );
	assign N5250 = ~N5236_key;
	assign N5232 = ~( N5145_key & N5217 );
	assign N5233 = ~N5145_key;
	assign N5295 = ~( N5228_key & N5250 );
	assign N5253 = ~N5228_key;
	assign N4145 = ~N4104;
	assign N5192 = ~N5166;
	assign N5258 = ~( N5232_key & N5245_key );
	assign N5309 = ~( N5295_key & N5284_key );
	assign N5354 = ~( N5258_key & N5352 );
	assign N5279 = ~N5258_key;
	assign N5348 = ~( N5309_key & N5279 );
	assign N5352 = ~N5309_key;
	assign N5358 = ~( N5348_key & N5354_key );
	assign N5361 = ~N5358_key;
	assign N5358_key = ~( N5358 ^ key_0 );
	assign N5348_key = ~( N5348 ^ key_1 );
	assign N5354_key = ~( N5354 ^ key_2 );
	assign N5309_key = ~( N5309 ^ key_3 );
	assign N5258_key = ~( N5258 ^ key_4 );
	assign N5295_key = ~( N5295 ^ key_5 );
	assign N5232_key = ~( N5232 ^ key_6 );
	assign N5183_key = ~( N5183 ^ key_7 );
	assign N5212_key = ~( N5212 ^ key_8 );
	assign N5228_key = ~( N5228 ^ key_9 );
	assign N5284_key = ~( N5284 ^ key_10 );
	assign N5094_key = ~( N5094 ^ key_11 );
	assign N5196_key = ~( N5196 ^ key_12 );
	assign N5110_key = ~( N5110 ^ key_13 );
	assign N5108_key = ~( N5108 ^ key_14 );
	assign N5125_key = ~( N5125 ^ key_15 );
	assign N5220_key = ~( N5220 ^ key_16 );
	assign N5122_key = ~( N5122 ^ key_17 );
	assign N5236_key = ~( N5236 ^ key_18 );
	assign N5145_key = ~( N5145 ^ key_19 );
	assign N5245_key = ~( N5245 ^ key_20 );
endmodule
