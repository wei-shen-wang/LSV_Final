module c3540(N343, N330, N326, N322, N317, N311, N303, N283, N274, N270, N257, N264, N250, N238, N68, N349, N223, N97, N20, N107, N13, N244, N41, N33, N294, N128, N116, N159, N350, N213, N45, N200, N77, N87, N143, N232, N58, N226, N1, N125, N132, N137, N150, N169, N329, N124, N179, N190, N50, N222, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, N5360, N5231, N5192, N5102, N5078, N5047, N1713, N5120, N4944, N1947, N3833, N5361, N5121, N4815, N3195, N4028, N3987, N4145, N5045, N4589, N4667, N5002);
	input N343, N330, N326, N322, N317, N311, N303, N283, N274, N270, N257, N264, N250, N238, N68, N349, N223, N97, N20, N107, N13, N244, N41, N33, N294, N128, N116, N159, N350, N213, N45, N200, N77, N87, N143, N232, N58, N226, N1, N125, N132, N137, N150, N169, N329, N124, N179, N190, N50, N222;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20;
	output N5360, N5231, N5192, N5102, N5078, N5047, N1713, N5120, N4944, N1947, N3833, N5361, N5121, N4815, N3195, N4028, N3987, N4145, N5045, N4589, N4667, N5002;
	wire N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350, N1562, N2482, N1325, N1667, N913, N1331, N914, N1756, N1821, N1761, N769, N1197, N1219, N1409, N793, N1452, N1337, N786, N890, N892, N1581, N1586, N1589, N1592, N1597, N1600, N2486, N2487, N794, N1117, N829, N2022, N2024, N2026, N2028, N2030, N2032, N2034, N2036, N1738, N1818, N820, N896, n_88, n_101, n_114, n_127, n_140, n_153, n_177, N832, N835, N1322, N3387, N3389, N1315, N839, N1520, N1792, N3216, N3225, N3234, N3243, N3252, N3261, N3270, N2068, N2348, N1251, N2133, N1870, N665, N1787, N1794, N3224, N3233, N3242, N3251, N3260, N3269, N2073, N2148, N1252, N1960, N1875, N679, N1729, N1789, N1796, N3232, N3241, N3250, N3259, N3268, N2078, N1253, N1267, N1727, N2134, N1880, N686, N1791, N1798, N3240, N3249, N3258, N3267, N2083, N1254, N2135, N1885, N702, N1714, N1793, N1800, N3248, N3257, N3266, N3275, N2088, N1255, N2136, N1890, N724, N1795, N1802, N3256, N3265, N3276, N3283, N3290, N2093, N1256, N1961, N2137, N1895, N736, N1797, N3264, N3277, N3284, N3291, N3298, N3305, N2098, N1257, N1730, N2138, N1900, N749, N1799, N2349, N3278, N3285, N3292, N3299, N3306, N3313, N3320, N2103, N1258, N2139, N1905, N763, N3207, N3214, N3215, N3213, N3222, N3223, N3212, N3221, N3230, N3231, N3211, N3220, N3229, N3238, N3239, N3210, N3219, N3228, N3237, N3246, N3247, N1788, N3209, N3218, N3227, N3236, N3245, N3254, N3255, N1790, N3208, N3217, N3226, N3235, N3244, N3253, N3262, N3263, N3407, N3423, N3431, N3439, N3455, N3463, N3645, N3664, N1179, N3410, N3426, N3434, N3442, N3458, N3466, N3648, N3667, n_73, N3383, N3413, N3429, N3437, N3445, N3461, N3469, N3651, N3670, N1358, N1803, N3414, N3430, N3438, N3446, N3462, N3470, N3652, N3671, N889, N1909, N5215, N1913, N920, N1643, N1644, N2023, N1645, N2025, N2417, N1510, N1259, N1646, N2027, N2420, N1509, N1260, N1647, N2029, N2425, N1512, N1261, N1648, N2031, N2430, N1511, N1262, N1067, N1649, N2033, N2435, N1692, N1467, N1650, N2035, N2438, N1691, N1468, N768, N2037, N2443, N1694, N1469, N2448, N1693, N1470, N2418, N2436, N2439, N1801, N3271, N3286, N3293, N3300, N3307, N3314, N3321, N3328, N3279, N3294, N3301, N3308, N3315, N3322, N3329, N3287, N3302, N3309, N3316, N3323, N3330, N3295, N3310, N3317, N3324, N3331, N3303, N3318, N3325, N3332, N3311, N3326, N3333, N3319, N3334, N3327, N4186, N4242, N4387, N4493, N4549, N4772, N4331, N4545, N4608, N4515, N1460, N4390, N4435, N1464, N2307, N2730, N2121, N2761, N1983, N1747, N1328, N2419, N2422, N2427, N2432, N2437, N2440, N2445, N2450, N2043, N1202, N2184, N1770, N2181, N2180, N2633, N2641, N2632, N2481, N1306, N4498, N1869, N1196, N1833, N1824, N1809, N891, N1806, N1366, N1986, N1987, N1988, N1989, N1990, N1991, N2768, N2769, N1580, N1579, N1426, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2144, N2143, N2211, n_164, N1850, N1815, n_83, n_96, n_109, n_122, n_135, n_148, n_172, N1401, N3552, N3544, N3546, N3550, N3548, N3540, N3542, N1893, N3534, N3536, N1898, N1966, N2350, N2376, N2758, n_145, n_169, n_94, n_107, n_134, n_121, n_79, N2652, N2478, N1507, N2325, N2398, N2898, N1250, N1940, n_161, n_93, n_133, n_82, N3419, N2146, N2899, N1263, n_150, n_106, n_120, N2666, N2328, N2900, n_174, n_132, n_162, n_81, N2677, N2901, N1505, N1947, n_98, n_119, n_151, N2688, N1508, N2331, N2347, N1340, n_111, n_80, n_163, n_175, N3451, N2147, N2351, N1264, n_137, n_152, n_99, N2706, N2334, N2355, N2483, n_176, n_112, n_124, N2719, N1722, N2353, n_157, n_160, n_159, n_144, n_147, n_168, n_158, n_171, n_92, n_146, n_95, n_105, n_170, n_108, n_131, n_118, N3644, N3657, N3661, N3663, N3676, N3680, N3789, N3803, n_74, N3471, N3557, N3568, N3573, N3578, N3589, N3594, N3731, N3753, N2185, N2188, N2197, N2200, N1353, N2206, N3172, N3682, N1912, N5231, N3175, N3178, N3181, N3184, N3187, N3605, N3690, N1917, N2656, N1715, N2659, N2670, N1718, N2681, N2692, N1933, N2697, N2710, N1936, N2723, n_149, n_100, n_138, n_85, n_173, n_113, n_125, n_97, n_139, n_86, n_110, n_126, n_136, n_87, n_123, n_84, N4675, N4291, N4678, N4461, N4786, N4596, N4716, N4558, N4924, N4706, N4859, N4817, N4468, N4589, N4644, N4559, N4463, N4788, N4602, N4708, N4507, N5136, N1461, N5277, N5286, N2310, N4350, N4341, N4344, N4347, N4475, N4472, N4335, N4338, N4647, N4794, N4800, N4831, N4838, N4907, N4913, N4985, N4588, N3195, N2145, N1673, N4921, N2764, N2379, N3406, N3642, N3779, N3780, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N4650, N4797, N4954, N4957, N4973, N5010, N5013, N5030, N1873, N2230, N2234, N2194, N1812, N2203, N2270, N2277, N2282, N2287, N2294, N2299, N3119, N3149, N2980, N3388, N3632, N3633, N3538, N3551, N3543, N3545, N3549, N3547, N3539, N3541, N3641, N3637, N3638, N3640, N3639, N3635, N3636, N2648, N1721, N2755, N2474, N3634, n_156, N1338, N3415, N2374, n_143, N2662, N2754, N2475, n_167, N2673, n_91, N1713, N2352, N2684, N2757, N2476, N3206, N1343, N3447, N2375, N3535, N2702, N2756, N2477, N3712, N4965, N2715, N1725, N3711, N3537, N3721, N3992, N3734, N3654, N3740, N3658, N3743, N3996, N3756, N3673, N3762, N3677, N3838, N3786, N3845, N3800, N3194, N2984, N2985, N2988, N2989, N2191, N2991, N4075, N3681, N4147, N3898, N3912, N4076, N3685, N4077, N3687, N4078, N3689, N4079, N3693, N4080, N3694, N4094, N4151, N3906, N3809, N3812, N3815, N3818, N3916, N4056, N4091, N3115, N2749, N2467, N3125, N3131, N2748, N2468, N3138, N3145, N2342, N2141, N3155, N3161, N2341, N2142, N3168, N4711, N4636, N4717, N4641, N4818, N4748, N4757, N4677, N4946, N4897, N4895, N4860, N4808, N4901, N4900, N4442, N4916, N4982, N4981, N4870, N4823, N4754, N4743, N4674, N5193, N5114, N5128, N5298, N5278, N5285, N4730, N4880, N4991, N4999, N5021, N5055, N5085, N5061, N4667, N2354, n_104, n_130, n_117, n_78, n_154, n_141, n_165, n_89, n_102, n_128, n_115, n_76, N4189, N4191, N4192, N4303, N4193, N4195, N4196, N4304, N2987, N2990, N2973, N2977, N5002, N3926, N3894, N4029, N3930, N3931, N4042, N4074, N4310, N4030, N4043, N4031, N4046, N3932, N3895, N4032, N3935, N3936, N4049, N4073, N4033, N4050, N4034, N4051, N4106, N4113, N4110, N4122, N2986, N4105, N4190, N3947, N4107, N4108, N4109, N4111, N4112, N4284, N4317, N4443, N4194, N4446, N3920, N4325, N4447, N4421, N4327, N4287, N4238, N4393, N4328, N4013, N3948, N4283, N4322, N4528, N4326, N4448, N4295, N2966, n_75, N2471, N4775, N4889, N4905, N4904, N4968, N4930, N4872, N4926, N4829, N4950, N4951, N5007, N4928, N4868, N4969, N4902, N5242, N5201, N5223, N5222, N5340, N5344, N5066, N5094, N4815, N5133, N5196, N4944, N5110, N5045, N5108, N5047, N5125, N5078, N5183, N5102, N5212, N5120, N5220, N5121, n_155, n_166, n_90, n_142, n_103, n_116, n_77, n_129, N3834, N3628, N3775, N3776, N4028, N4104, N4733, N4562, N4705, N4146, N4572, N4252, N4503, N4552, N4148, N4487, N4149, N4555, N4150, N4319, N4329, N4152, N4153, N4668, N4506, N4629, N4630, N4573, N4256, N4416, N4509, N4508, N4427, N4530, N4496, N4458, N4576, N3706, N3196, N3705, N3627, N4953, N4906, N4983, N4970, N5254, N5360, N5350, N5166, N5122, N5236, N5145, N5228, N3987, N4145, N4769, N4688, N4740, N4670, N4619, N4527, N4669, N4593, N4599, N4511, N4704, N4623, N4526, N4510, N4640, N4635, N3773, N4931, N4984, N5266, N5192, N5245, N5217, N5284, N5250, N5232, N5233, N5295, N5253, N4816, N4896, N4673, N4747, N4753, N4676, N3833, N5258, N5309, N5354, N5279, N5348, N5352, N5358, N5361;
	wire N5358_key, N5348_key, N5354_key, N5309_key, N5258_key, N5183_key, N5212_key, N5228_key, N5284_key, N5295_key, N5094_key, N5196_key, N5110_key, N5108_key, N5125_key, N5220_key, N5122_key, N5236_key, N5145_key, N5245_key, N5232_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20;
	assign N1562 = ( N1 & N1337 );
	assign N2482 = ( N1761 & N1 );
	assign N1325 = ( N1 & N786 & N20 );
	assign N1667 = ( N1 & N13 & N1426 );
	assign N913 = ~( N1 & N13 );
	assign N1331 = ~( N1 & N786 );
	assign N914 = ~( N1 & N20 & N33 );
	assign N1756 = ~( N1 & N13 & N20 );
	assign N1821 = ~( N1 & N13 & N1179 );
	assign N1761 = ~( N1 & N786 & N20 & N832 );
	assign N769 = ~N1;
	assign N1197 = ( N794 | N1 );
	assign N1219 = ( N820 | N1 );
	assign N1409 = ( N1 | N1196 );
	assign N793 = ( N13 & N20 );
	assign N1452 = ( N769 & N13 & N794 );
	assign N1337 = ~( N13 & N794 & N45 );
	assign N786 = ~N13;
	assign N890 = ( N20 & N200 );
	assign N892 = ( N20 & N179 );
	assign N1581 = ( N1338 & N20 );
	assign N1586 = ( N686 & N20 );
	assign N1589 = ( N77 & N20 );
	assign N1592 = ( N1343 & N20 );
	assign N1597 = ( N749 & N20 );
	assign N1600 = ( N116 & N20 );
	assign N2486 = ( N2374 & N20 );
	assign N2487 = ( N2375 & N20 );
	assign N794 = ~N20;
	assign N1117 = ( N820 | N20 );
	assign N829 = ( N33 & N41 );
	assign N2022 = ( N77 & N33 );
	assign N2024 = ( N87 & N33 );
	assign N2026 = ( N97 & N33 );
	assign N2028 = ( N107 & N33 );
	assign N2030 = ( N116 & N33 );
	assign N2032 = ( N283 & N33 );
	assign N2034 = ( N294 & N33 );
	assign N2036 = ( N303 & N33 );
	assign N1738 = ~( N1325 & N33 );
	assign N1818 = ~( N33 & N832 );
	assign N820 = ~N33;
	assign N896 = ( N349 | N33 );
	assign n_88 = ( n_84 & N33 );
	assign n_101 = ( n_97 & N33 );
	assign n_114 = ( n_110 & N33 );
	assign n_127 = ( n_123 & N33 );
	assign n_140 = ( n_136 & N33 );
	assign n_153 = ( n_149 & N33 );
	assign n_177 = ( n_173 & N33 );
	assign N832 = ~N41;
	assign N835 = ( N41 | N45 );
	assign N1322 = ( N769 & N45 );
	assign N3387 = ( N3196 & N45 );
	assign N3389 = ( N2973 & N45 );
	assign N1315 = ( N769 & N45 & N832 );
	assign N839 = ~N45;
	assign N1520 = ( N50 & N1263 );
	assign N1792 = ( N50 & N1580 );
	assign N3216 = ( N50 & N2985 );
	assign N3225 = ( N50 & N2986 );
	assign N3234 = ( N50 & N2987 );
	assign N3243 = ( N50 & N2988 );
	assign N3252 = ( N50 & N2989 );
	assign N3261 = ( N50 & N2990 );
	assign N3270 = ( N50 & N2991 );
	assign N2068 = ( N50 & N1197 & N1869 );
	assign N2348 = ( N2146 & N77 & N50 );
	assign N1251 = ~( N226 & N50 );
	assign N2133 = ~( N50 & N58 );
	assign N1870 = ~( N50 | N1409 );
	assign N665 = ~N50;
	assign N1787 = ( N58 & N1579 );
	assign N1794 = ( N58 & N1580 );
	assign N3224 = ( N58 & N2985 );
	assign N3233 = ( N58 & N2986 );
	assign N3242 = ( N58 & N2987 );
	assign N3251 = ( N58 & N2988 );
	assign N3260 = ( N58 & N2989 );
	assign N3269 = ( N58 & N2990 );
	assign N2073 = ( N58 & N1197 & N1869 );
	assign N2148 = ( N1722 & N1267 & N665 & N58 );
	assign N1252 = ~( N232 & N58 );
	assign N1960 = ~( N58 & N686 );
	assign N1875 = ~( N58 | N1409 );
	assign N679 = ~N58;
	assign N1729 = ( N68 & N665 );
	assign N1789 = ( N68 & N1579 );
	assign N1796 = ( N68 & N1580 );
	assign N3232 = ( N68 & N2985 );
	assign N3241 = ( N68 & N2986 );
	assign N3250 = ( N68 & N2987 );
	assign N3259 = ( N68 & N2988 );
	assign N3268 = ( N68 & N2989 );
	assign N2078 = ( N68 & N1197 & N1869 );
	assign N1253 = ~( N238 & N68 );
	assign N1267 = ~( N68 & N77 );
	assign N1727 = ~( N68 & N679 );
	assign N2134 = ~( N702 & N68 );
	assign N1880 = ~( N68 | N1409 );
	assign N686 = ~N68;
	assign N1791 = ( N77 & N1579 );
	assign N1798 = ( N77 & N1580 );
	assign N3240 = ( N77 & N2985 );
	assign N3249 = ( N77 & N2986 );
	assign N3258 = ( N77 & N2987 );
	assign N3267 = ( N77 & N2988 );
	assign N2083 = ( N77 & N1197 & N1869 );
	assign N1254 = ~( N244 & N77 );
	assign N2135 = ~( N686 & N77 );
	assign N1885 = ~( N77 | N1409 );
	assign N702 = ~N77;
	assign N1714 = ( N87 & N1264 );
	assign N1793 = ( N87 & N1579 );
	assign N1800 = ( N87 & N1580 );
	assign N3248 = ( N87 & N2985 );
	assign N3257 = ( N87 & N2986 );
	assign N3266 = ( N87 & N2987 );
	assign N3275 = ( N87 & N2988 );
	assign N2088 = ( N87 & N1219 & N1869 );
	assign N1255 = ~( N250 & N87 );
	assign N2136 = ~( N736 & N87 );
	assign N1890 = ~( N87 | N1409 );
	assign N724 = ~N87;
	assign N1795 = ( N97 & N1579 );
	assign N1802 = ( N97 & N1580 );
	assign N3256 = ( N97 & N2985 );
	assign N3265 = ( N97 & N2986 );
	assign N3276 = ( N97 & N2989 );
	assign N3283 = ( N97 & N2988 );
	assign N3290 = ( N97 & N2987 );
	assign N2093 = ( N97 & N1219 & N1869 );
	assign N1256 = ~( N257 & N97 );
	assign N1961 = ~( N97 & N749 );
	assign N2137 = ~( N724 & N97 );
	assign N1895 = ~( N97 | N1409 );
	assign N736 = ~N97;
	assign N1797 = ( N107 & N1579 );
	assign N3264 = ( N107 & N2985 );
	assign N3277 = ( N107 & N2990 );
	assign N3284 = ( N107 & N2989 );
	assign N3291 = ( N107 & N2988 );
	assign N3298 = ( N107 & N2987 );
	assign N3305 = ( N107 & N2986 );
	assign N2098 = ( N107 & N1219 & N1869 );
	assign N1257 = ~( N264 & N107 );
	assign N1730 = ~( N107 & N736 );
	assign N2138 = ~( N763 & N107 );
	assign N1900 = ~( N107 | N1409 );
	assign N749 = ~N107;
	assign N1799 = ( N116 & N1579 );
	assign N2349 = ( N116 & N2147 );
	assign N3278 = ( N116 & N2991 );
	assign N3285 = ( N116 & N2990 );
	assign N3292 = ( N116 & N2989 );
	assign N3299 = ( N116 & N2988 );
	assign N3306 = ( N116 & N2987 );
	assign N3313 = ( N116 & N2986 );
	assign N3320 = ( N116 & N2985 );
	assign N2103 = ( N116 & N1219 & N1869 );
	assign N1258 = ~( N270 & N116 );
	assign N2139 = ~( N749 & N116 );
	assign N1905 = ~( N116 | N1409 );
	assign N763 = ~N116;
	assign N3207 = ( N124 & N2984 );
	assign N3214 = ( N125 & N2991 );
	assign N3215 = ( N125 & N2984 );
	assign N3213 = ( N128 & N2990 );
	assign N3222 = ( N128 & N2991 );
	assign N3223 = ( N128 & N2984 );
	assign N3212 = ( N132 & N2989 );
	assign N3221 = ( N132 & N2990 );
	assign N3230 = ( N132 & N2991 );
	assign N3231 = ( N132 & N2984 );
	assign N3211 = ( N137 & N2988 );
	assign N3220 = ( N137 & N2989 );
	assign N3229 = ( N137 & N2990 );
	assign N3238 = ( N137 & N2991 );
	assign N3239 = ( N137 & N2984 );
	assign N3210 = ( N143 & N2987 );
	assign N3219 = ( N143 & N2988 );
	assign N3228 = ( N143 & N2989 );
	assign N3237 = ( N143 & N2990 );
	assign N3246 = ( N143 & N2991 );
	assign N3247 = ( N143 & N2984 );
	assign N1788 = ( N150 & N1580 );
	assign N3209 = ( N150 & N2986 );
	assign N3218 = ( N150 & N2987 );
	assign N3227 = ( N150 & N2988 );
	assign N3236 = ( N150 & N2989 );
	assign N3245 = ( N150 & N2990 );
	assign N3254 = ( N150 & N2991 );
	assign N3255 = ( N150 & N2984 );
	assign N1790 = ( N159 & N1580 );
	assign N3208 = ( N159 & N2985 );
	assign N3217 = ( N159 & N2986 );
	assign N3226 = ( N159 & N2987 );
	assign N3235 = ( N159 & N2988 );
	assign N3244 = ( N159 & N2989 );
	assign N3253 = ( N159 & N2990 );
	assign N3262 = ( N159 & N2991 );
	assign N3263 = ( N159 & N2984 );
	assign N3407 = ( N169 & N2648 & N2656 );
	assign N3423 = ( N169 & N2662 & N2670 );
	assign N3431 = ( N169 & N2673 & N2681 );
	assign N3439 = ( N169 & N2684 & N2692 );
	assign N3455 = ( N169 & N2702 & N2710 );
	assign N3463 = ( N169 & N2715 & N2723 );
	assign N3645 = ( N169 & N3415 & N2659 );
	assign N3664 = ( N169 & N3447 & N2697 );
	assign N1179 = ( N794 | N169 );
	assign N3410 = ( N179 & N2648 & N3115 );
	assign N3426 = ( N179 & N2662 & N3131 );
	assign N3434 = ( N179 & N2673 & N3138 );
	assign N3442 = ( N179 & N2684 & N3145 );
	assign N3458 = ( N179 & N2702 & N3161 );
	assign N3466 = ( N179 & N2715 & N3168 );
	assign N3648 = ( N179 & N3415 & N3125 );
	assign N3667 = ( N179 & N3447 & N3155 );
	assign n_73 = ~N179;
	assign N3383 = ( N3161 & N3168 & N179 & n_75 );
	assign N3413 = ( N190 & N2652 & N3115 );
	assign N3429 = ( N190 & N2666 & N3131 );
	assign N3437 = ( N190 & N2677 & N3138 );
	assign N3445 = ( N190 & N2688 & N3145 );
	assign N3461 = ( N190 & N2706 & N3161 );
	assign N3469 = ( N190 & N2719 & N3168 );
	assign N3651 = ( N190 & N3419 & N3125 );
	assign N3670 = ( N190 & N3451 & N3155 );
	assign N1358 = ~( N794 | N190 );
	assign N1803 = ( N200 & N892 );
	assign N3414 = ( N200 & N2652 & N2656 );
	assign N3430 = ( N200 & N2666 & N2670 );
	assign N3438 = ( N200 & N2677 & N2681 );
	assign N3446 = ( N200 & N2688 & N2692 );
	assign N3462 = ( N200 & N2706 & N2710 );
	assign N3470 = ( N200 & N2719 & N2723 );
	assign N3652 = ( N200 & N3419 & N2659 );
	assign N3671 = ( N200 & N3451 & N2697 );
	assign N889 = ~N200;
	assign N1909 = ( N1452 & N213 );
	assign N5215 = ( N213 & N5193 );
	assign N1913 = ( N1452 & N213 & N343 );
	assign N920 = ~N213;
	assign N1643 = ( N222 & N1401 );
	assign N1644 = ( N223 & N1401 );
	assign N2023 = ( N223 & N1850 );
	assign N1645 = ( N226 & N1401 );
	assign N2025 = ( N226 & N1850 );
	assign N2417 = ( N2043 & N226 & N1873 );
	assign N1510 = ~( N226 & N1260 );
	assign N1259 = ~N226;
	assign N1646 = ( N232 & N1401 );
	assign N2027 = ( N232 & N1850 );
	assign N2420 = ( N2043 & N232 & N1873 );
	assign N1509 = ~( N232 & N1259 );
	assign N1260 = ~N232;
	assign N1647 = ( N238 & N1401 );
	assign N2029 = ( N238 & N1850 );
	assign N2425 = ( N2043 & N238 & N1873 );
	assign N1512 = ~( N238 & N1262 );
	assign N1261 = ~N238;
	assign N1648 = ( N244 & N1401 );
	assign N2031 = ( N244 & N1850 );
	assign N2430 = ( N2043 & N244 & N1873 );
	assign N1511 = ~( N244 & N1261 );
	assign N1262 = ~N244;
	assign N1067 = ( N250 & N768 );
	assign N1649 = ( N250 & N1401 );
	assign N2033 = ( N250 & N1850 );
	assign N2435 = ( N2043 & N250 & N1893 );
	assign N1692 = ~( N250 & N1468 );
	assign N1467 = ~N250;
	assign N1650 = ( N257 & N1401 );
	assign N2035 = ( N257 & N1850 );
	assign N2438 = ( N2043 & N257 & N1898 );
	assign N1691 = ~( N257 & N1467 );
	assign N1468 = ~N257;
	assign N768 = ( N257 | N264 );
	assign N2037 = ( N264 & N1850 );
	assign N2443 = ( N2043 & N264 & N1898 );
	assign N1694 = ~( N264 & N1470 );
	assign N1469 = ~N264;
	assign N2448 = ( N2043 & N270 & N1898 );
	assign N1693 = ~( N270 & N1469 );
	assign N1470 = ~N270;
	assign N2418 = ( N2043 & N274 & N1306 );
	assign N2436 = ( N2043 & N274 & N1322 );
	assign N2439 = ( N2043 & N274 & N1315 );
	assign N1801 = ( N283 & N1579 );
	assign N3271 = ( N283 & N2984 );
	assign N3286 = ( N283 & N2991 );
	assign N3293 = ( N283 & N2990 );
	assign N3300 = ( N283 & N2989 );
	assign N3307 = ( N283 & N2988 );
	assign N3314 = ( N283 & N2987 );
	assign N3321 = ( N283 & N2986 );
	assign N3328 = ( N283 & N2985 );
	assign N3279 = ( N294 & N2984 );
	assign N3294 = ( N294 & N2991 );
	assign N3301 = ( N294 & N2990 );
	assign N3308 = ( N294 & N2989 );
	assign N3315 = ( N294 & N2988 );
	assign N3322 = ( N294 & N2987 );
	assign N3329 = ( N294 & N2986 );
	assign N3287 = ( N303 & N2984 );
	assign N3302 = ( N303 & N2991 );
	assign N3309 = ( N303 & N2990 );
	assign N3316 = ( N303 & N2989 );
	assign N3323 = ( N303 & N2988 );
	assign N3330 = ( N303 & N2987 );
	assign N3295 = ( N311 & N2984 );
	assign N3310 = ( N311 & N2991 );
	assign N3317 = ( N311 & N2990 );
	assign N3324 = ( N311 & N2989 );
	assign N3331 = ( N311 & N2988 );
	assign N3303 = ( N317 & N2984 );
	assign N3318 = ( N317 & N2991 );
	assign N3325 = ( N317 & N2990 );
	assign N3332 = ( N317 & N2989 );
	assign N3311 = ( N322 & N2984 );
	assign N3326 = ( N322 & N2991 );
	assign N3333 = ( N322 & N2990 );
	assign N3319 = ( N326 & N2984 );
	assign N3334 = ( N326 & N2991 );
	assign N3327 = ( N329 & N2984 );
	assign N4186 = ( N330 & N4094 );
	assign N4242 = ( N330 & N4112 );
	assign N4387 = ( N330 & N4317 );
	assign N4493 = ( N330 & N4319 );
	assign N4549 = ( N330 & N4443 );
	assign N4772 = ( N330 & N4704 );
	assign N4331 = ( N330 & N4094 & N4295 );
	assign N4545 = ( N330 & N4319 & N4496 );
	assign N4608 = ( N330 & N4284 & N4562 );
	assign N4515 = ~( N330 & N4153 );
	assign N1460 = ~N330;
	assign N4390 = ( N330 & N4112 & N4111 & N4194 );
	assign N4435 = ( N330 & N4094 & N4108 & N4107 );
	assign N1464 = ~( N920 | N343 );
	assign N2307 = ( N1464 & N350 );
	assign N2730 = ( N1562 & N1761 );
	assign N2121 = ~N1562;
	assign N2761 = ( N1722 & N2482 );
	assign N1983 = ( N1067 & N1325 );
	assign N1747 = ~( N1325 & N820 );
	assign N1328 = ~N1325;
	assign N2419 = ( N1667 & N2238 );
	assign N2422 = ( N1667 & N2239 );
	assign N2427 = ( N1667 & N2240 );
	assign N2432 = ( N1667 & N2241 );
	assign N2437 = ( N1667 & N2242 );
	assign N2440 = ( N1667 & N2243 );
	assign N2445 = ( N1667 & N2244 );
	assign N2450 = ( N1667 & N2245 );
	assign N2043 = ~N1667;
	assign N1202 = ( N913 & N914 );
	assign N2184 = ( N1331 & N1756 );
	assign N1770 = ~N1331;
	assign N2181 = ( N1756 & N1328 );
	assign N2180 = ~N1756;
	assign N2633 = ( N1821 & N1833 );
	assign N2641 = ( N1821 & N1824 );
	assign N2632 = ~N1821;
	assign N2481 = ~N1761;
	assign N1306 = ( N769 & N835 );
	assign N4498 = ( N4442 & N769 );
	assign N1869 = ( N1202 & N1409 );
	assign N1196 = ~N793;
	assign N1833 = ~( N786 & N820 );
	assign N1824 = ~( N786 & N794 & N820 );
	assign N1809 = ( N890 & N1366 );
	assign N891 = ~N890;
	assign N1806 = ( N889 & N892 );
	assign N1366 = ~N892;
	assign N1986 = ( N1581 | N1787 | N1788 );
	assign N1987 = ( N1586 | N1791 | N1792 );
	assign N1988 = ( N1589 | N1793 | N1794 );
	assign N1989 = ( N1592 | N1795 | N1796 );
	assign N1990 = ( N1597 | N1799 | N1800 );
	assign N1991 = ( N1600 | N1801 | N1802 );
	assign N2768 = ( N2486 | N1789 | N1790 );
	assign N2769 = ( N2487 | N1797 | N1798 );
	assign N1580 = ( N794 & N1117 );
	assign N1579 = ~N1117;
	assign N1426 = ~N829;
	assign N2238 = ( N2022 | N1643 | N2023 );
	assign N2239 = ( N2024 | N1644 | N2025 );
	assign N2240 = ( N2026 | N1645 | N2027 );
	assign N2241 = ( N2028 | N1646 | N2029 );
	assign N2242 = ( N2030 | N1647 | N2031 );
	assign N2243 = ( N2032 | N1648 | N2033 );
	assign N2244 = ( N2034 | N1649 | N2035 );
	assign N2245 = ( N2036 | N1650 | N2037 );
	assign N2144 = ( N1738 & N1747 );
	assign N2143 = ~N1738;
	assign N2211 = ( N1815 & N1818 );
	assign n_164 = ~( N3278 | N1818 );
	assign N1850 = ( N820 & N896 );
	assign N1815 = ~( N820 & N832 );
	assign n_83 = ( n_79 & N820 );
	assign n_96 = ( n_92 & N820 );
	assign n_109 = ( n_105 & N820 );
	assign n_122 = ( n_118 & N820 );
	assign n_135 = ( n_131 & N820 );
	assign n_148 = ( n_144 & N820 );
	assign n_172 = ( n_168 & N820 );
	assign N1401 = ~N896;
	assign N3552 = ( n_85 & n_86 & n_87 & n_88 );
	assign N3544 = ( n_98 & n_99 & n_100 & n_101 );
	assign N3546 = ( n_111 & n_112 & n_113 & n_114 );
	assign N3550 = ( n_124 & n_125 & n_126 & n_127 );
	assign N3548 = ( n_137 & n_138 & n_139 & n_140 );
	assign N3540 = ( n_150 & n_151 & n_152 & n_153 );
	assign N3542 = ( n_174 & n_175 & n_176 & n_177 );
	assign N1893 = ~N1322;
	assign N3534 = ~( N3387 | N2350 );
	assign N3536 = ~( N3389 | N1966 );
	assign N1898 = ~N1315;
	assign N1966 = ( N1520 & N839 );
	assign N2350 = ( N2148 & N839 );
	assign N2376 = ( N1520 & N2180 );
	assign N2758 = ( N1520 & N2481 );
	assign n_145 = ~( N3215 | N3216 | N3217 );
	assign n_169 = ~( N3223 | N3224 | N3225 );
	assign n_94 = ~( N3234 | N3235 );
	assign n_107 = ~( N3242 | N3243 );
	assign n_134 = ~( N3252 | N3253 );
	assign n_121 = ~( N3260 | N3261 );
	assign n_79 = ~N3270;
	assign N2652 = ~( N2270 | N1870 | N2068 );
	assign N2478 = ( N2348 | N1729 );
	assign N1507 = ( N1251 & N1252 & N1253 & N1254 );
	assign N2325 = ~( N1940 & N2133 );
	assign N2398 = ( N665 & N2211 );
	assign N2898 = ( N665 & N2633 );
	assign N1250 = ( N665 & N679 & N686 );
	assign N1940 = ~( N679 & N665 );
	assign n_161 = ~( N3271 | N3224 | N3241 );
	assign n_93 = ~( N3231 | N3232 | N3233 );
	assign n_133 = ~( N3250 | N3251 );
	assign n_82 = ~( N3268 | N3269 );
	assign N3419 = ~( N3119 | N1875 | N2073 );
	assign N2146 = ~( N1727 & N1960 );
	assign N2899 = ( N679 & N2633 );
	assign N1263 = ~( N679 & N686 );
	assign n_150 = ~( N3279 | N3232 | N3249 );
	assign n_106 = ~( N3239 | N3240 | N3241 );
	assign n_120 = ~( N3258 | N3259 );
	assign N2666 = ~( N2277 | N1880 | N2078 );
	assign N2328 = ~( N2134 & N2135 );
	assign N2900 = ( N686 & N2633 );
	assign n_174 = ~( N3287 | N3240 | N3257 );
	assign n_132 = ~( N3247 | N3248 | N3249 );
	assign n_162 = ~( N3258 | N3275 );
	assign n_81 = ~( N3266 | N3267 );
	assign N2677 = ~( N2282 | N1885 | N2083 );
	assign N2901 = ( N702 & N2633 );
	assign N1505 = ~( N702 & N1250 );
	assign N1947 = ~N1714;
	assign n_98 = ~( N3295 | N3248 | N3265 );
	assign n_119 = ~( N3255 | N3256 | N3257 );
	assign n_151 = ~( N3266 | N3283 );
	assign N2688 = ~( N2287 | N1890 | N2088 );
	assign N1508 = ( N1255 & N1256 & N1257 & N1258 );
	assign N2331 = ~( N2136 & N2137 );
	assign N2347 = ( N724 & N2144 );
	assign N1340 = ( N724 & N736 & N749 );
	assign n_111 = ~( N3303 | N3256 | N3305 );
	assign n_80 = ~( N3263 | N3264 | N3265 );
	assign n_163 = ~( N3276 | N3277 );
	assign n_175 = ~( N3290 | N3291 );
	assign N3451 = ~( N3149 | N1895 | N2093 );
	assign N2147 = ~( N1730 & N1961 );
	assign N2351 = ( N736 & N2144 );
	assign N1264 = ~( N736 & N749 );
	assign n_137 = ~( N3311 | N3264 | N3313 );
	assign n_152 = ~( N3284 | N3285 );
	assign n_99 = ~( N3298 | N3299 );
	assign N2706 = ~( N2294 | N1900 | N2098 );
	assign N2334 = ~( N2138 & N2139 );
	assign N2355 = ( N749 & N2144 );
	assign N2483 = ( N2349 & N2180 );
	assign n_176 = ~( N3292 | N3293 );
	assign n_112 = ~( N3306 | N3307 );
	assign n_124 = ~( N3319 | N3320 | N3321 );
	assign N2719 = ~( N2299 | N1905 | N2103 );
	assign N1722 = ( N763 & N1340 );
	assign N2353 = ( N763 & N2144 );
	assign n_157 = ~( N3207 | N3208 | N3209 );
	assign n_160 = ~( N3214 | N1815 );
	assign n_159 = ~( N3212 | N3213 );
	assign n_144 = ~N3222;
	assign n_147 = ~( N3220 | N3221 );
	assign n_168 = ~N3230;
	assign n_158 = ~( N3210 | N3211 );
	assign n_171 = ~( N3228 | N3229 );
	assign n_92 = ~N3238;
	assign n_146 = ~( N3218 | N3219 );
	assign n_95 = ~( N3236 | N3237 );
	assign n_105 = ~N3246;
	assign n_170 = ~( N3226 | N3227 );
	assign n_108 = ~( N3244 | N3245 );
	assign n_131 = ~N3254;
	assign n_118 = ~N3262;
	assign N3644 = ~( N3407 | N3410 );
	assign N3657 = ~( N3423 | N3426 );
	assign N3661 = ~( N3431 | N3434 );
	assign N3663 = ~( N3439 | N3442 );
	assign N3676 = ~( N3455 | N3458 );
	assign N3680 = ~( N3463 | N3466 );
	assign N3789 = ~( N3645 | N3648 );
	assign N3803 = ~( N3664 | N3667 );
	assign n_74 = ( n_73 & N2692 );
	assign N3471 = ( N3194 | N3383 );
	assign N3557 = ( N3413 | N3414 | N2648 );
	assign N3568 = ( N3429 | N3430 | N2662 );
	assign N3573 = ( N3437 | N3438 | N2673 );
	assign N3578 = ( N3445 | N3446 | N2684 );
	assign N3589 = ( N3461 | N3462 | N2702 );
	assign N3594 = ( N3469 | N3470 | N2715 );
	assign N3731 = ( N3651 | N3652 | N3415 );
	assign N3753 = ( N3670 | N3671 | N3447 );
	assign N2185 = ~( N1358 & N1812 );
	assign N2188 = ~( N1358 & N1809 );
	assign N2197 = ~( N1358 & N1806 );
	assign N2200 = ~( N1358 & N1803 );
	assign N1353 = ~N1358;
	assign N2206 = ~( N1353 & N1803 );
	assign N3172 = ( N1909 & N2648 );
	assign N3682 = ( N1909 & N3415 );
	assign N1912 = ~N1909;
	assign N5231 = ~N5215;
	assign N3175 = ( N1913 & N2662 );
	assign N3178 = ( N1913 & N2673 );
	assign N3181 = ( N1913 & N2684 );
	assign N3184 = ( N1913 & N2702 );
	assign N3187 = ( N1913 & N2715 );
	assign N3605 = ( N3471 & N1913 );
	assign N3690 = ( N1913 & N3447 );
	assign N1917 = ~N1913;
	assign N2656 = ( N2417 | N2418 | N2419 );
	assign N1715 = ~( N1509 & N1510 );
	assign N2659 = ( N2420 | N2418 | N2422 );
	assign N2670 = ( N2425 | N2418 | N2427 );
	assign N1718 = ~( N1511 & N1512 );
	assign N2681 = ( N2430 | N2418 | N2432 );
	assign N2692 = ( N2435 | N2436 | N2437 );
	assign N1933 = ~( N1691 & N1692 );
	assign N2697 = ( N2438 | N2439 | N2440 );
	assign N2710 = ( N2443 | N2439 | N2445 );
	assign N1936 = ~( N1693 & N1694 );
	assign N2723 = ( N2448 | N2439 | N2450 );
	assign n_149 = ~N3286;
	assign n_100 = ~( N3300 | N3301 );
	assign n_138 = ~( N3314 | N3315 );
	assign n_85 = ~( N3327 | N3328 | N3329 );
	assign n_173 = ~N3294;
	assign n_113 = ~( N3308 | N3309 );
	assign n_125 = ~( N3322 | N3323 );
	assign n_97 = ~N3302;
	assign n_139 = ~( N3316 | N3317 );
	assign n_86 = ~( N3330 | N3331 );
	assign n_110 = ~N3310;
	assign n_126 = ~( N3324 | N3325 );
	assign n_136 = ~N3318;
	assign n_87 = ~( N3332 | N3333 );
	assign n_123 = ~N3326;
	assign n_84 = ~N3334;
	assign N4675 = ~( N4186 & N4635 );
	assign N4291 = ~N4186;
	assign N4678 = ~( N4242 & N4640 );
	assign N4461 = ~N4242;
	assign N4786 = ~( N4387 & N4747 );
	assign N4596 = ~N4387;
	assign N4716 = ~( N4493 & N4676 );
	assign N4558 = ~N4493;
	assign N4924 = ~( N4549 & N4896 );
	assign N4706 = ~N4549;
	assign N4859 = ~( N4772 & N4816 );
	assign N4817 = ~N4772;
	assign N4468 = ~( N4331 | N4091 );
	assign N4589 = ( N4545 | N4287 );
	assign N4644 = ~( N4608 | N4310 );
	assign N4559 = ~( N4463 & N4515 );
	assign N4463 = ~( N4112 & N1460 );
	assign N4788 = ~( N4390 & N4753 );
	assign N4602 = ~N4390;
	assign N4708 = ~( N4435 & N4673 );
	assign N4507 = ~N4435;
	assign N5136 = ( N5055 & N5085 & N1464 );
	assign N1461 = ~N1464;
	assign N5277 = ( N5236_key & N5254 & N2307 );
	assign N5286 = ( N5250 & N5266 & N2307 );
	assign N2310 = ~N2307;
	assign N4350 = ( n_76 & n_77 & n_78 & N2730 );
	assign N4341 = ( n_89 & n_90 & n_91 & N2730 );
	assign N4344 = ( n_102 & n_103 & n_104 & N2730 );
	assign N4347 = ( n_115 & n_116 & n_117 & N2730 );
	assign N4475 = ( n_128 & n_129 & n_130 & N2730 );
	assign N4472 = ( n_141 & n_142 & n_143 & N2730 );
	assign N4335 = ( n_154 & n_155 & n_156 & N2730 );
	assign N4338 = ( n_165 & n_166 & n_167 & N2730 );
	assign N4647 = ( N4559 & N2121 );
	assign N4794 = ( N4711 & N2121 );
	assign N4800 = ( N4717 & N2121 );
	assign N4831 = ( N4743 & N2121 );
	assign N4838 = ( N4757 & N2121 );
	assign N4907 = ( N4818 & N2121 );
	assign N4913 = ( N4823 & N2121 );
	assign N4985 = ( N4946 & N2121 );
	assign N4588 = ~( N2758 | N4498 | N2761 );
	assign N3195 = ~( N2376 | N1983 | N2379 );
	assign N2145 = ~N1747;
	assign N1673 = ~N1202;
	assign N4921 = ( N4895 & N2184 );
	assign N2764 = ( N2478 & N1770 );
	assign N2379 = ( N1721 & N2181 );
	assign N3406 = ( N3206 & N2641 );
	assign N3642 = ( N3535 & N2641 );
	assign N3779 = ( N3712 & N2641 );
	assign N3780 = ( N3711 & N2641 );
	assign N3713 = ( N3634 & N2632 );
	assign N3714 = ( N3635 & N2632 );
	assign N3715 = ( N3636 & N2632 );
	assign N3716 = ( N3637 & N2632 );
	assign N3717 = ( N3638 & N2632 );
	assign N3718 = ( N3639 & N2632 );
	assign N3719 = ( N3640 & N2632 );
	assign N3720 = ( N3641 & N2632 );
	assign N4650 = ( N4559 & N2481 );
	assign N4797 = ( N4711 & N2481 );
	assign N4954 = ( N4926 & N2481 );
	assign N4957 = ( N4931 & N2481 );
	assign N4973 = ( N4953 & N2481 );
	assign N5010 = ( N4983 & N2481 );
	assign N5013 = ( N4984 & N2481 );
	assign N5030 = ( N5007 & N2481 );
	assign N1873 = ~N1306;
	assign N2230 = ~N1833;
	assign N2234 = ~N1824;
	assign N2194 = ~( N1353 & N1809 );
	assign N1812 = ( N891 & N1366 );
	assign N2203 = ~( N1353 & N1806 );
	assign N2270 = ( N1986 & N1673 );
	assign N2277 = ( N1987 & N1673 );
	assign N2282 = ( N1988 & N1673 );
	assign N2287 = ( N1989 & N1673 );
	assign N2294 = ( N1990 & N1673 );
	assign N2299 = ( N1991 & N1673 );
	assign N3119 = ( N2768 & N1673 );
	assign N3149 = ( N2769 & N1673 );
	assign N2980 = ( N2471 & N2143 );
	assign N3388 = ( N2977 & N2143 );
	assign N3632 = ( N3536 & N2143 );
	assign N3633 = ( N3534 & N2143 );
	assign N3538 = ( n_161 & n_162 & n_163 & n_164 );
	assign N3551 = ( n_80 & n_81 & n_82 & n_83 );
	assign N3543 = ( n_93 & n_94 & n_95 & n_96 );
	assign N3545 = ( n_106 & n_107 & n_108 & n_109 );
	assign N3549 = ( n_119 & n_120 & n_121 & n_122 );
	assign N3547 = ( n_132 & n_133 & n_134 & n_135 );
	assign N3539 = ( n_145 & n_146 & n_147 & n_148 );
	assign N3541 = ( n_169 & n_170 & n_171 & n_172 );
	assign N3641 = ( N3551 | N3552 );
	assign N3637 = ( N3543 | N3544 );
	assign N3638 = ( N3545 | N3546 );
	assign N3640 = ( N3549 | N3550 );
	assign N3639 = ( N3547 | N3548 );
	assign N3635 = ( N3539 | N3540 );
	assign N3636 = ( N3541 | N3542 );
	assign N2648 = ~N2652;
	assign N1721 = ~( N1507 & N1508 );
	assign N2755 = ~( N2325 & N2475 );
	assign N2474 = ~N2325;
	assign N3634 = ( N3537 | N3538 | N2398 );
	assign n_156 = ~N2898;
	assign N1338 = ~N1250;
	assign N3415 = ~N3419;
	assign N2374 = ~N2146;
	assign n_143 = ~N2899;
	assign N2662 = ~N2666;
	assign N2754 = ~( N2328 & N2474 );
	assign N2475 = ~N2328;
	assign n_167 = ~N2900;
	assign N2673 = ~N2677;
	assign n_91 = ~N2901;
	assign N1713 = ~N1505;
	assign N2352 = ( N1947 & N2145 );
	assign N2684 = ~N2688;
	assign N2757 = ~( N2331 & N2477 );
	assign N2476 = ~N2331;
	assign N3206 = ( N2980 | N2145 | N2347 );
	assign N1343 = ~N1340;
	assign N3447 = ~N3451;
	assign N2375 = ~N2147;
	assign N3535 = ( N3388 | N2145 | N2351 );
	assign N2702 = ~N2706;
	assign N2756 = ~( N2334 & N2476 );
	assign N2477 = ~N2334;
	assign N3712 = ( N3633 | N2354 | N2355 );
	assign N4965 = ~( N2764 | N2483 | N4921 );
	assign N2715 = ~N2719;
	assign N1725 = ~N1722;
	assign N3711 = ( N3632 | N2352 | N2353 );
	assign N3537 = ( n_157 & n_158 & n_159 & n_160 );
	assign N3721 = ( N3644 & N3557 );
	assign N3992 = ~( N3644 & N3894 & N3930 & N3931 );
	assign N3734 = ( N3657 & N3568 );
	assign N3654 = ~N3657;
	assign N3740 = ( N3661 & N3573 );
	assign N3658 = ~N3661;
	assign N3743 = ( N3663 & N3578 );
	assign N3996 = ~( N3663 & N3895 & N3935 & N3936 );
	assign N3756 = ( N3676 & N3589 );
	assign N3673 = ~N3676;
	assign N3762 = ( N3680 & N3594 );
	assign N3677 = ~N3680;
	assign N3838 = ( N3789 & N3731 );
	assign N3786 = ~N3789;
	assign N3845 = ( N3803 & N3753 );
	assign N3800 = ~N3803;
	assign N3194 = ( N2697 & N2710 & N2723 & n_74 );
	assign N2984 = ~N2185;
	assign N2985 = ~N2188;
	assign N2988 = ~N2197;
	assign N2989 = ~N2200;
	assign N2191 = ~( N1353 & N1812 );
	assign N2991 = ~N2206;
	assign N4075 = ~( N3172 & N4042 );
	assign N3681 = ~N3172;
	assign N4147 = ~( N3682 & N4113 );
	assign N3898 = ~N3682;
	assign N3912 = ( N3786 & N1912 );
	assign N4076 = ~( N3175 & N4043 );
	assign N3685 = ~N3175;
	assign N4077 = ~( N3178 & N4046 );
	assign N3687 = ~N3178;
	assign N4078 = ~( N3181 & N4049 );
	assign N3689 = ~N3181;
	assign N4079 = ~( N3184 & N4050 );
	assign N3693 = ~N3184;
	assign N4080 = ~( N3187 & N4051 );
	assign N3694 = ~N3187;
	assign N4094 = ( N3605 | N4056 );
	assign N4151 = ~( N3690 & N4122 );
	assign N3906 = ~N3690;
	assign N3809 = ( N3654 & N1917 );
	assign N3812 = ( N3658 & N1917 );
	assign N3815 = ( N3673 & N1917 );
	assign N3818 = ( N3677 & N1917 );
	assign N3916 = ( N3800 & N1917 );
	assign N4056 = ( N3932 & N1917 );
	assign N4091 = ( N3996 & N1917 );
	assign N3115 = ~N2656;
	assign N2749 = ~( N1715 & N2468 );
	assign N2467 = ~N1715;
	assign N3125 = ~N2659;
	assign N3131 = ~N2670;
	assign N2748 = ~( N1718 & N2467 );
	assign N2468 = ~N1718;
	assign N3138 = ~N2681;
	assign N3145 = ~N2692;
	assign N2342 = ~( N1933 & N2142 );
	assign N2141 = ~N1933;
	assign N3155 = ~N2697;
	assign N3161 = ~N2710;
	assign N2341 = ~( N1936 & N2141 );
	assign N2142 = ~N1936;
	assign N3168 = ~N2723;
	assign N4711 = ~( N4675 & N4636 );
	assign N4636 = ~( N4576 & N4291 );
	assign N4717 = ~( N4678 & N4641 );
	assign N4641 = ~( N4458 & N4461 );
	assign N4818 = ~( N4786 & N4748 );
	assign N4748 = ~( N4593 & N4596 );
	assign N4757 = ~( N4716 & N4677 );
	assign N4677 = ~( N4623 & N4558 );
	assign N4946 = ~( N4924 & N4897 );
	assign N4897 = ~( N4740 & N4706 );
	assign N4895 = ~( N4859 & N4860 );
	assign N4860 = ~( N4769 & N4817 );
	assign N4808 = ( N4717 & N4468 );
	assign N4901 = ( N4717 & N4757 & N4823 & N4468 );
	assign N4900 = ~( N4868 | N4468 );
	assign N4442 = ~N4468;
	assign N4916 = ( N4818 & N4644 );
	assign N4982 = ( N4818 & N4743 & N4946 & N4644 );
	assign N4981 = ~( N4968 | N4644 );
	assign N4870 = ~N4644;
	assign N4823 = ~( N4788 & N4754 );
	assign N4754 = ~( N4599 & N4602 );
	assign N4743 = ~( N4708 & N4674 );
	assign N4674 = ~( N4619 & N4507 );
	assign N5193 = ~( N5136 | N5166 );
	assign N5114 = ( N5102 & N1461 );
	assign N5128 = ( N1461 & N5120 );
	assign N5298 = ( N5277 | N5285 | N5278 | N5286 );
	assign N5278 = ( N5250 & N5254 & N2310 );
	assign N5285 = ( N5236_key & N5266 & N2310 );
	assign N4730 = ~( N4647 | N4650 | N4350 );
	assign N4880 = ~( N4794 | N4797 | N4341 );
	assign N4991 = ~( N4913 | N4954 | N4344 );
	assign N4999 = ~( N4800 | N4957 | N4347 );
	assign N5021 = ~( N4838 | N4973 | N4475 );
	assign N5055 = ~( N4831 | N5010 | N4472 );
	assign N5085 = ~( N4985 | N5030 | N4335 );
	assign N5061 = ~( N4907 | N5013 | N4338 );
	assign N4667 = ~N4588;
	assign N2354 = ( N1725 & N2145 );
	assign n_104 = ~N3406;
	assign n_130 = ~N3642;
	assign n_117 = ~N3779;
	assign n_78 = ~N3780;
	assign n_154 = ~N3713;
	assign n_141 = ~N3714;
	assign n_165 = ~N3715;
	assign n_89 = ~N3716;
	assign n_102 = ~N3717;
	assign n_128 = ~N3718;
	assign n_115 = ~N3719;
	assign n_76 = ~N3720;
	assign N4189 = ( N4146 & N2230 );
	assign N4191 = ( N4148 & N2230 );
	assign N4192 = ( N4149 & N2230 );
	assign N4303 = ( N4252 & N2230 );
	assign N4193 = ( N4150 & N2234 );
	assign N4195 = ( N4152 & N2234 );
	assign N4196 = ( N4153 & N2234 );
	assign N4304 = ( N4256 & N2234 );
	assign N2987 = ~N2194;
	assign N2990 = ~N2203;
	assign N2973 = ~( N2754 & N2755 );
	assign N2977 = ~( N2756 & N2757 );
	assign N5002 = ~N4965;
	assign N3926 = ( N3721 & N3838 & N3734 & N3740 );
	assign N3894 = ~( N3721 & N3786 );
	assign N4029 = ~( N3721 & N3681 );
	assign N3930 = ~( N3721 & N3838 & N3654 );
	assign N3931 = ~( N3658 & N3838 & N3734 & N3721 );
	assign N4042 = ~N3721;
	assign N4074 = ~N3992;
	assign N4310 = ( N3992 | N4283 );
	assign N4030 = ~( N3734 & N3685 );
	assign N4043 = ~N3734;
	assign N4031 = ~( N3740 & N3687 );
	assign N4046 = ~N3740;
	assign N3932 = ( N3743 & N3845 & N3756 & N3762 );
	assign N3895 = ~( N3743 & N3800 );
	assign N4032 = ~( N3743 & N3689 );
	assign N3935 = ~( N3743 & N3845 & N3673 );
	assign N3936 = ~( N3677 & N3845 & N3756 & N3743 );
	assign N4049 = ~N3743;
	assign N4073 = ~( N3926 & N3996 );
	assign N4033 = ~( N3756 & N3693 );
	assign N4050 = ~N3756;
	assign N4034 = ~( N3762 & N3694 );
	assign N4051 = ~N3762;
	assign N4106 = ~( N3838 & N3898 );
	assign N4113 = ~N3838;
	assign N4110 = ~( N3845 & N3906 );
	assign N4122 = ~N3845;
	assign N2986 = ~N2191;
	assign N4105 = ~( N4075 & N4029 );
	assign N4190 = ~( N4147 & N4106 );
	assign N3947 = ~N3912;
	assign N4107 = ~( N4076 & N4030 );
	assign N4108 = ~( N4077 & N4031 );
	assign N4109 = ~( N4078 & N4032 );
	assign N4111 = ~( N4079 & N4033 );
	assign N4112 = ~( N4080 & N4034 );
	assign N4284 = ( N4094 & N3926 );
	assign N4317 = ( N4094 & N4108 );
	assign N4443 = ( N4094 & N4190 & N4107 & N4108 );
	assign N4194 = ~( N4151 & N4110 );
	assign N4446 = ~( N4190 & N3809 );
	assign N3920 = ~N3809;
	assign N4325 = ~( N4107 & N3812 );
	assign N4447 = ~( N4190 & N4107 & N3812 );
	assign N4421 = ( N3812 | N4322 );
	assign N4327 = ~( N4194 & N3815 );
	assign N4287 = ( N3815 | N4238 );
	assign N4238 = ( N4111 & N3818 );
	assign N4393 = ~( N3818 & N4152 );
	assign N4328 = ~( N4194 & N4111 & N3818 );
	assign N4013 = ~N3818;
	assign N3948 = ~N3916;
	assign N4283 = ( N4091 & N3926 );
	assign N4322 = ( N4091 & N4108 );
	assign N4528 = ~( N4091 & N4149 );
	assign N4326 = ~( N4107 & N4108 & N4091 );
	assign N4448 = ~( N4190 & N4107 & N4108 & N4091 );
	assign N4295 = ~N4091;
	assign N2966 = ~( N2748 & N2749 );
	assign n_75 = ( N3145 & N3155 );
	assign N2471 = ~( N2341 & N2342 );
	assign N4775 = ~N4717;
	assign N4889 = ~N4818;
	assign N4905 = ~( N4757 & N4872 );
	assign N4904 = ~N4757;
	assign N4968 = ~N4946;
	assign N4930 = ~( N4808 & N4904 );
	assign N4872 = ~N4808;
	assign N4926 = ( N4900 | N4901 );
	assign N4829 = ~( N4775 & N4442 );
	assign N4950 = ~( N4916 & N4902 );
	assign N4951 = ~N4916;
	assign N5007 = ( N4981 | N4982 );
	assign N4928 = ~( N4889 & N4870 );
	assign N4868 = ~N4823;
	assign N4969 = ~( N4743 & N4951 );
	assign N4902 = ~N4743;
	assign N5242 = ~( N5114 & N5222 );
	assign N5201 = ~N5114;
	assign N5223 = ~( N5128 & N5201 );
	assign N5222 = ~N5128;
	assign N5340 = ~( N5298 & N5258_key );
	assign N5344 = ~N5298;
	assign N5066 = ( N4730 & N4999 & N5021 & N4991 );
	assign N5094 = ~( N5047 & N4730 );
	assign N4815 = ~N4730;
	assign N5133 = ( N4880 & N5061 & N5055 & N5085 );
	assign N5196 = ~( N5121 & N4880 );
	assign N4944 = ~N4880;
	assign N5110 = ~( N5078 & N4991 );
	assign N5045 = ~N4991;
	assign N5108 = ~( N4815 & N4999 );
	assign N5047 = ~N4999;
	assign N5125 = ~( N5045 & N5021 );
	assign N5078 = ~N5021;
	assign N5183 = ~( N5120 & N5055 );
	assign N5102 = ~N5055;
	assign N5212 = ~( N5102 & N5085 );
	assign N5120 = ~N5085;
	assign N5220 = ~( N4944 & N5061 );
	assign N5121 = ~N5061;
	assign n_155 = ~N4189;
	assign n_166 = ~N4191;
	assign n_90 = ~N4192;
	assign n_142 = ~N4303;
	assign n_103 = ~N4193;
	assign n_116 = ~N4195;
	assign n_77 = ~N4196;
	assign n_129 = ~N4304;
	assign N3834 = ~( N2973 & N3776 );
	assign N3628 = ~N2973;
	assign N3775 = ~( N2977 & N3628 );
	assign N3776 = ~N2977;
	assign N4028 = ( N3932 & N3926 );
	assign N4104 = ( N4073 & N4074 );
	assign N4733 = ~( N4310 & N4669 );
	assign N4562 = ~N4310;
	assign N4705 = ~( N4105 & N4669 );
	assign N4146 = ~N4105;
	assign N4572 = ~( N4190 & N4526 );
	assign N4252 = ~N4190;
	assign N4503 = ~( N3947 & N4446 & N4447 & N4448 );
	assign N4552 = ~( N4107 & N4508 );
	assign N4148 = ~N4107;
	assign N4487 = ~( N4108 & N4295 );
	assign N4149 = ~N4108;
	assign N4555 = ~( N4109 & N4510 );
	assign N4150 = ~N4109;
	assign N4319 = ( N4112 & N4111 );
	assign N4329 = ~( N4111 & N4013 );
	assign N4152 = ~N4111;
	assign N4153 = ~N4112;
	assign N4668 = ~( N4284 & N4630 );
	assign N4506 = ~N4284;
	assign N4629 = ~( N4443 & N4506 );
	assign N4630 = ~N4443;
	assign N4573 = ~( N4194 & N4496 );
	assign N4256 = ~N4194;
	assign N4416 = ~( N3920 & N4325 & N4326 );
	assign N4509 = ~( N4421 & N4148 );
	assign N4508 = ~N4421;
	assign N4427 = ~( N3948 & N4327 & N4328 );
	assign N4530 = ~( N4287 & N4256 );
	assign N4496 = ~N4287;
	assign N4458 = ~( N4329 & N4393 );
	assign N4576 = ~( N4487 & N4528 );
	assign N3706 = ~( N2966 & N3627 );
	assign N3196 = ~N2966;
	assign N3705 = ~( N2471 & N3196 );
	assign N3627 = ~N2471;
	assign N4953 = ~( N4930 & N4905 );
	assign N4906 = ~( N4872 & N4829 );
	assign N4983 = ~( N4950 & N4969 );
	assign N4970 = ~( N4951 & N4928 );
	assign N5254 = ~( N5242 & N5223 );
	assign N5360 = ~( N5350 & N5340 );
	assign N5350 = ~( N5279 & N5344 );
	assign N5166 = ( N5066 & N5133 );
	assign N5122 = ~( N5094_key & N5108_key );
	assign N5236 = ~( N5196_key & N5220_key );
	assign N5145 = ~( N5125_key & N5110_key );
	assign N5228 = ~( N5183_key & N5212_key );
	assign N3987 = ~( N3775 & N3834 );
	assign N4145 = ~N4104;
	assign N4769 = ~( N4733 & N4688 );
	assign N4688 = ~( N4503 & N4562 );
	assign N4740 = ~( N4705 & N4670 );
	assign N4670 = ~( N4503 & N4146 );
	assign N4619 = ~( N4572 & N4527 );
	assign N4527 = ~( N4416 & N4252 );
	assign N4669 = ~N4503;
	assign N4593 = ~( N4552 & N4509 );
	assign N4599 = ~( N4555 & N4511 );
	assign N4511 = ~( N4427 & N4150 );
	assign N4704 = ~( N4629 & N4668 );
	assign N4623 = ~( N4573 & N4530 );
	assign N4526 = ~N4416;
	assign N4510 = ~N4427;
	assign N4640 = ~N4458;
	assign N4635 = ~N4576;
	assign N3773 = ~( N3705 & N3706 );
	assign N4931 = ~N4906;
	assign N4984 = ~N4970;
	assign N5266 = ~N5254;
	assign N5192 = ~N5166;
	assign N5245 = ~( N5122_key & N5233 );
	assign N5217 = ~N5122_key;
	assign N5284 = ~( N5236_key & N5253 );
	assign N5250 = ~N5236_key;
	assign N5232 = ~( N5145_key & N5217 );
	assign N5233 = ~N5145_key;
	assign N5295 = ~( N5228_key & N5250 );
	assign N5253 = ~N5228_key;
	assign N4816 = ~N4769;
	assign N4896 = ~N4740;
	assign N4673 = ~N4619;
	assign N4747 = ~N4593;
	assign N4753 = ~N4599;
	assign N4676 = ~N4623;
	assign N3833 = ~N3773;
	assign N5258 = ~( N5232_key & N5245_key );
	assign N5309 = ~( N5295_key & N5284_key );
	assign N5354 = ~( N5258_key & N5352 );
	assign N5279 = ~N5258_key;
	assign N5348 = ~( N5309_key & N5279 );
	assign N5352 = ~N5309_key;
	assign N5358 = ~( N5348_key & N5354_key );
	assign N5361 = ~N5358_key;
	assign N5358_key = ~( N5358 ^ key_0 );
	assign N5348_key = ~( N5348 ^ key_1 );
	assign N5354_key = ~( N5354 ^ key_2 );
	assign N5309_key = ~( N5309 ^ key_3 );
	assign N5258_key = ~( N5258 ^ key_4 );
	assign N5183_key = ~( N5183 ^ key_5 );
	assign N5212_key = ~( N5212 ^ key_6 );
	assign N5228_key = ~( N5228 ^ key_7 );
	assign N5284_key = ~( N5284 ^ key_8 );
	assign N5295_key = ~( N5295 ^ key_9 );
	assign N5094_key = ~( N5094 ^ key_10 );
	assign N5196_key = ~( N5196 ^ key_11 );
	assign N5110_key = ~( N5110 ^ key_12 );
	assign N5108_key = ~( N5108 ^ key_13 );
	assign N5125_key = ~( N5125 ^ key_14 );
	assign N5220_key = ~( N5220 ^ key_15 );
	assign N5122_key = ~( N5122 ^ key_16 );
	assign N5236_key = ~( N5236 ^ key_17 );
	assign N5145_key = ~( N5145 ^ key_18 );
	assign N5245_key = ~( N5245 ^ key_19 );
	assign N5232_key = ~( N5232 ^ key_20 );
endmodule
