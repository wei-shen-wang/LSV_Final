module c5315(N1, N100, N103, N106, N109, N11, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N14, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N17, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N20, N200, N203, N206, N209, N210, N217, N218, N225, N226, N23, N233, N234, N24, N241, N242, N245, N248, N25, N251, N254, N257, N26, N264, N265, N27, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N31, N315, N316, N323, N324, N331, N332, N335, N338, N34, N341, N348, N351, N358, N361, N366, N369, N37, N372, N373, N374, N386, N389, N4, N40, N400, N411, N422, N43, N435, N446, N457, N46, N468, N479, N49, N490, N503, N514, N52, N523, N53, N534, N54, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N61, N610, N613, N616, N619, N625, N631, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N709, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474_key, N7476_key, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128, N816);
	input N1, N100, N103, N106, N109, N11, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N14, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N17, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N20, N200, N203, N206, N209, N210, N217, N218, N225, N226, N23, N233, N234, N24, N241, N242, N245, N248, N25, N251, N254, N257, N26, N264, N265, N27, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N31, N315, N316, N323, N324, N331, N332, N335, N338, N34, N341, N348, N351, N358, N361, N366, N369, N37, N372, N373, N374, N386, N389, N4, N40, N400, N411, N422, N43, N435, N446, N457, N46, N468, N479, N49, N490, N503, N514, N52, N523, N53, N534, N54, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N61, N610, N613, N616, N619, N625, N631, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123;
	output N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N709, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474_key, N7476_key, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128, N816;
	wire N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, N3360, N3359, N3358, N3357, N2309, N1146, N6107, N6664, AND3_1351_inw1, AND4_1349_inw1, N6806, N2637, AND3_600_inw1, AND3_619_inw1, AND3_609_inw1, AND3_617_inw1, AND3_230_inw1, AND3_238_inw1, AND3_229_inw1, AND3_237_inw1, AND3_813_inw1, AND3_807_inw1, AND3_808_inw1, AND3_809_inw1, N1150, N1475, N3740, AND3_228_inw1, AND3_236_inw1, AND3_227_inw1, AND3_235_inw1, AND3_605_inw1, AND3_613_inw1, AND3_602_inw1, AND3_610_inw1, AND3_225_inw1, AND3_233_inw1, AND3_733_inw1, AND3_730_inw1, N5119, N6693, AND3_1400_inw1, AND4_1398_inw1, N5955, N2715, AND3_223_inw1, AND3_244_inw1, AND3_232_inw1, AND3_240_inw1, AND3_608_inw1, AND3_616_inw1, AND3_231_inw1, AND3_239_inw1, AND3_607_inw1, AND3_615_inw1, AND3_606_inw1, AND3_614_inw1, AND3_812_inw1, AND3_815_inw1, AND3_810_inw1, AND3_814_inw1, N2969, N3738, N2970, N3739, N2971, AND3_604_inw1, AND3_612_inw1, N3072, N3071, AND3_603_inw1, AND3_611_inw1, AND3_226_inw1, AND3_234_inw1, AND3_222_inw1, AND3_224_inw1, AND3_597_inw1, AND3_601_inw1, AND3_734_inw1, AND3_729_inw1, AND3_731_inw1, AND3_732_inw1, AND3_735_inw1, AND3_717_inw1, AND3_620_inw1, AND3_723_inw1, AND3_618_inw1, AND3_736_inw1, AND3_728_inw1, AND3_242_inw1, AND3_737_inw1, AND3_718_inw1, AND3_719_inw1, AND3_720_inw1, AND3_722_inw1, AND3_724_inw1, AND3_721_inw1, N6880, N6478, N1042, N2054, N2139, N7506, N7511, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8125, N8126, N2590, N2142, N709, N1147, N4737, N4738, N4739, N4740, AND3_212_inw1, AND3_221_inw1, AND3_583_inw1, AND3_594_inw1, AND3_211_inw1, AND3_220_inw1, AND3_582_inw1, AND3_593_inw1, AND3_210_inw1, AND3_219_inw1, AND3_207_inw1, AND3_217_inw1, AND3_206_inw1, AND3_216_inw1, AND3_205_inw1, AND3_215_inw1, AND3_203_inw1, AND3_213_inw1, AND3_204_inw1, AND3_214_inw1, AND3_621_inw1, AND3_622_inw1, AND3_271_inw1, AND3_292_inw1, AND3_580_inw1, AND3_591_inw1, AND3_209_inw1, AND3_218_inw1, AND3_581_inw1, AND3_592_inw1, AND3_579_inw1, AND3_590_inw1, AND3_578_inw1, AND3_589_inw1, AND3_577_inw1, AND3_588_inw1, AND3_575_inw1, AND3_586_inw1, AND3_576_inw1, AND3_587_inw1, N3689, N3761, N3758, N3823, N3753, N2876, N2835, N3027, N3688, N2831, N3023, N4024, N2823, N2875, N2836, N3028, N3687, N2832, N3024, N3610, N2825, N2874, N2837, N3029, N3686, N2833, N3025, N3609, N2827, N2873, N2838, N3030, N3685, N2834, N3026, N3563, N2829, N2872, N2910, N2911, N2912, N2938, N2939, N2940, N2941, N2983, N2985, N2986, N2984, N1152, n_331, N2907, N2980, N3013, AND3_351_inw1, AND3_352_inw1, AND3_377_inw1, AND3_378_inw1, AND3_379_inw1, AND3_380_inw1, AND3_408_inw1, AND3_410_inw1, AND3_411_inw1, AND3_444_inw1, AND3_445_inw1, AND3_446_inw1, AND3_447_inw1, AND3_700_inw1, N3444, N3502, AND3_512_inw1, AND3_513_inw1, AND3_524_inw1, AND3_525_inw1, AND3_526_inw1, AND3_527_inw1, AND3_532_inw1, AND3_534_inw1, AND3_535_inw1, AND3_547_inw1, AND3_548_inw1, AND3_549_inw1, AND3_550_inw1, AND3_790_inw1, N3447, N3448, N3449, N3463, N3464, N3465, N3466, N3485, N3486, N3487, N3508, N3509, N3510, N3511, N3982, N2851, N3684, N2847, N2934, N3562, N2839, N2871, N2852, N3683, N2848, N2935, N3561, N2841, N2870, N2853, N3682, N2849, N2936, N3560, N2843, N2869, N2854, N3681, N2850, N2937, N3559, N2845, N2868, N3680, N3558, N3142, N2867, N816, N3731, N3608, N2901, N3604, N2527, N2963, N3613, N3730, N3607, N2902, N2962, N3729, N2908, N3606, N2903, N2961, N3728, N2909, N3605, N2905, N2960, N2923, N3727, N2919, N2979, N4953, N4954, N1660, N2959, N2954, N2955, N2956, N2957, N2958, N2942, N2855, N1144, N2924, N3726, N2921, N2981, N3515, N2915, N1138, N2925, N3725, N2922, N2982, N3514, N2917, N1145, N3724, N3513, N2999, N1139, N3723, N3512, N3032, N4310, AND3_324_inw1, AND3_506_inw1, N5250, N4608, N2636, N3679, N3722, N1151, g45_inw1, N4298, AND3_321_inw1, AND3_503_inw1, N5247, N2633, N3676, N3719, N4301, AND3_322_inw1, AND3_504_inw1, N5248, N2634, N3677, N3720, N4305, AND3_323_inw1, AND3_505_inw1, N5249, N2635, N3678, N3721, N4290, AND3_307_inw1, AND3_497_inw1, N5245, N4575, N2631, N3670, N3769, N4297, AND3_308_inw1, AND3_498_inw1, N5246, N2632, N3671, N3770, N4268, N5242, N2628, N4185, N4280, AND3_305_inw1, AND3_495_inw1, N5243, N2629, N3668, N3767, N4284, AND3_306_inw1, AND3_496_inw1, N5244, N2630, N3669, N3768, N4379, N5261, N2709, N3703, N4385, N5262, N4627, N2710, N3704, N4392, AND3_362_inw1, AND3_517_inw1, N5263, N2711, N3711, N3745, N2349, N4067, N5112, N2712, N2350, N4396, AND3_364_inw1, AND3_518_inw1, N5274, N2713, N3712, N3746, N4400, AND3_365_inw1, AND3_519_inw1, N5275, N2714, N3713, N3747, N1137, N2387, N1141, N1140, N1153, n_330, N1155, n_329, N1154, N8041, N7990, N7991, N1157, AND3_1879_inw1, AND3_1915_inw1, AND3_1917_inw1, AND3_1919_inw1, AND3_1921_inw1, AND3_2034_inw1, AND3_2036_inw1, AND3_2038_inw1, AND3_2040_inw1, AND3_2297_inw1, N2653, N2585, N2586, N2587, N2588, N2589, N2591, N2592, N2593, N2594, N2703, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3662, N2664, AND3_1881_inw1, AND3_1923_inw1, AND3_1925_inw1, AND3_1927_inw1, AND3_1929_inw1, AND3_2042_inw1, AND3_2044_inw1, AND3_2046_inw1, AND3_2048_inw1, AND3_2299_inw1, N2728, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2778, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3663, N2739, N8035, N7996, N7997, N1219, N3615, N1588, N1043, N1066, N1148, N1067, N1080, N1092, N1104, N2624, N7464, N1755, AND3_1792_inw1, AND3_1945_inw1, N1758, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N2790, AND3_1883_inw1, AND3_1932_inw1, AND3_1934_inw1, AND3_1936_inw1, AND3_1937_inw1, AND3_2052_inw1, AND3_2054_inw1, AND3_2056_inw1, AND3_2058_inw1, AND3_2293_inw1, N2779, AND3_1887_inw1, AND3_1939_inw1, AND3_1941_inw1, AND3_1943_inw1, AND3_1944_inw1, AND3_2050_inw1, AND3_2060_inw1, AND3_2062_inw1, AND3_2064_inw1, AND3_2295_inw1, N2801, N2604, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2626, N3638, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3660, N2812, N2625, N8077, N8078, AND3_1589_inw1, AND3_1803_inw1, AND3_1804_inw1, AND3_1834_inw1, AND3_1835_inw1, AND3_1836_inw1, AND3_1838_inw1, AND3_1839_inw1, AND3_1844_inw1, AND3_1845_inw1, AND3_1958_inw1, AND3_1959_inw1, AND3_1960_inw1, AND3_1961_inw1, AND3_1962_inw1, AND3_1963_inw1, AND3_1964_inw1, AND3_1965_inw1, AND3_2274_inw1, AND3_2275_inw1, N3068, N3659, N3661, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3063, N1972, N6512, g32_inw2, N6817, N6106, N6104, N6932, N6650, N4038, N4032, N4033, N4034, N2060, N4031, N4036, N4042, N4035, N4037, N4039, N4040, N2623, N3829, N5346, g28_inw2, N6844, N6163, N6161, N6164, N5616, N3831, N3828, N8096, N8093, N6979, N6879, N1149, N8127, N8128, N3893, OR3_836_inw1, N4183, N4264, N3980, OR3_627_inw1, OR3_709_inw1, N3887, N3664, N3763, N3405, N3401, N3504, OR3_628_inw1, OR3_710_inw1, N3881, N3665, N3764, N3824, N3406, N3402, N3505, OR3_629_inw1, OR3_711_inw1, N3873, N3666, N3765, N3407, N3403, N3506, OR3_630_inw1, OR3_712_inw1, N3867, N3667, N3766, N3797, N3408, N3404, N3507, N3705, OR3_653_inw1, OR3_654_inw1, OR3_666_inw1, OR3_667_inw1, OR3_668_inw1, OR3_669_inw1, OR3_687_inw1, OR3_688_inw1, OR3_689_inw1, N3816, g49_inw2, N3700, N3482, N3757, N3445, N3446, N3459, N3460, N3461, N3462, N3481, N3483, N3484, OR3_635_inw1, N3861, N3672, N3715, N3413, N3409, OR3_636_inw1, N3855, N3673, N3716, N3793, N3414, N3410, OR3_637_inw1, N3849, N3674, N3717, N3415, N3411, OR3_638_inw1, N3842, N3675, N3718, N3789, N3416, N3412, N4011, N3968, N3810, N3962, N3956, N3701, N3813, N3948, N3702, OR3_659_inw1, N3942, N3708, N3742, N5147, N5148, N3453, N3450, N4196, N4955, N4008, N3921, N3927, N3933, N3732, OR3_660_inw1, N3709, N3743, N3775, N3454, N3451, OR3_661_inw1, N3710, N3744, N3455, N3452, N3771, N6105, N6103, AND4_1345_inw2, N6990, N5728, g12_inw1, N5462, N6987, N5176, N5086, N4109, N4198, N2061, N6094, NOR4_1525_inw1, n_316, N5431, N5080, N4100, N4234, N6098, N6095, NOR3_1524_inw1, OR4_1517_inw1, OR4_1522_inw1, N5441, N5082, N4103, N4225, N6102, AND3_1344_inw1, AND4_1341_inw2, N6419, OR3_1518_inw1, N5452, N5084, N4106, N4228, N6088, AND3_1331_inw1, AND4_1322_inw2, N6816, N7153, N5469, N5418, N6815, N7152, N5087, N5076, N4094, N4240, n_306, N5424, N5078, N4097, N4231, OR4_1486_inw1, N5389, N5070, N4939, N6071, NOR3_1513_inw1, OR4_1512_inw1, N5396, N5072, N4088, N4243, N6083, N6072, N6494, OR3_1514_inw1, N5407, N5074, N4091, N4237, N5117, N5066, N6575, OR3_1528_inw1, N5562, N5107, N4144, N6146, AND3_1382_inw1, AND4_1323_inw2, N6843, N7159, N5622, N5573, N6842, N7158, N5120, N5109, N4147, n_308, N5579, N5111, N4153, N4252, N2920, N6152, NOR4_1538_inw1, n_314, N5264, N4856, N3456, N5954, N6153, NOR3_1537_inw1, OR4_1531_inw1, OR4_1535_inw1, N5595, N5114, N4156, N4246, N6159, AND3_1393_inw1, AND4_1391_inw2, N6445, OR3_1532_inw1, N5606, N5116, N4159, N4249, N1143, N1142, N2584, g49_inw1, N8045, OR4_2241_inw2, N8043, N7988, N7989, N7338, N7434, N7436, N7438, N7440, N7667, N7669, N7671, N7673, N8118, AND3_1743_inw1, AND3_1880_inw1, AND3_1914_inw1, AND3_1918_inw1, AND3_1920_inw1, AND3_2033_inw1, AND3_2035_inw1, AND3_2037_inw1, AND3_2039_inw1, AND3_2296_inw1, OR4_1974_inw2, OR4_2088_inw2, OR4_2089_inw2, OR4_2090_inw2, OR4_2091_inw2, OR4_1916_inw2, OR4_1976_inw2, OR4_1977_inw2, OR4_1978_inw2, OR4_2300_inw2, N7011, N7339, N7433, N7437, N7439, N7666, N7668, N7670, N7672, N8117, N7340, N7442, N7444, N7446, N7448, N7675, N7677, N7679, N7681, N8120, AND3_1744_inw1, AND3_1882_inw1, AND3_1922_inw1, AND3_1926_inw1, AND3_1928_inw1, AND3_2041_inw1, AND3_2043_inw1, AND3_2045_inw1, AND3_2047_inw1, AND3_2298_inw1, OR4_1979_inw2, OR4_2092_inw2, OR4_2093_inw2, OR4_2094_inw2, OR4_2095_inw2, OR4_1924_inw2, OR4_1981_inw2, OR4_1982_inw2, OR4_1983_inw2, OR4_2301_inw2, N7012, N7341, N7441, N7445, N7447, N7674, N7676, N7678, N7680, N8119, N8048, OR4_2242_inw2, N8044, N7994, N7995, OR4_873_inw2, OR4_874_inw2, OR4_876_inw2, OR4_877_inw2, N3614, OR4_1992_inw2, N4741, N7114, AND3_995_inw1, OR4_1930_inw2, OR4_2097_inw2, OR4_2098_inw2, OR4_2099_inw2, OR4_2100_inw2, OR4_1984_inw2, OR4_1985_inw2, OR4_1986_inw2, OR4_1987_inw2, OR4_2302_inw2, N7013, N7342, N7349, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N8113, N8114, AND3_1745_inw1, AND3_1884_inw1, AND3_1931_inw1, AND3_1933_inw1, AND3_1935_inw1, AND3_2051_inw1, AND3_2053_inw1, AND3_2055_inw1, AND3_2057_inw1, AND3_2292_inw1, N7364, N7458, N7460, N7462, N7463, N7683, N7693, N7695, N7697, N8116, AND3_1747_inw1, AND3_1885_inw1, AND3_1938_inw1, AND3_1940_inw1, AND3_1942_inw1, AND3_2049_inw1, AND3_2059_inw1, AND3_2061_inw1, AND3_2063_inw1, AND3_2294_inw1, OR4_2096_inw2, OR4_2101_inw2, OR4_2102_inw2, OR4_2103_inw2, OR4_1988_inw2, OR4_1989_inw2, OR4_1990_inw2, OR4_1991_inw2, OR4_2303_inw2, OR4_1950_inw2, N7016, N7357, N7457, N7459, N7461, N7682, N7692, N7694, N7696, N8115, OR4_2278_inw2, OR4_2279_inw2, N8079, N8082, N6718, N7146, N7147, N7187, N7188, N7189, N7196, N7197, N7207, N7208, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N8071, N8072, N7479, N7530, AND3_800_inw1, AND3_841_inw1, AND3_923_inw1, AND3_1006_inw1, AND3_1007_inw1, AND3_1008_inw1, AND3_1009_inw1, AND3_1010_inw1, AND3_1011_inw1, AND3_1024_inw1, AND3_1025_inw1, AND3_1026_inw1, AND3_1027_inw1, AND3_1028_inw1, AND3_1029_inw1, AND3_1030_inw1, AND3_1031_inw1, AND3_1139_inw1, AND3_1993_inw1, AND3_2029_inw1, N7190, N7270, N7276, N7282, N6866, N7198, N7288, N7294, N7304, N7531, N7537, N7543, N7549, N7310, N7555, N7561, N7567, N7573, N8089, N8090, N3998, N4197, N4547, N4956, N4957, N4958, N4959, N4960, N4961, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5165, N7526, N7636, N6830, N6829, N6101, N7040, N7125, N7126, N7127, N7023, N6508, OR4_1517_inw2, g33_inw1, OR4_876_inw1, OR4_873_inw1, OR4_874_inw1, N4272, N4275, N4279, OR4_877_inw1, N6856, N5956, N6158, N7064, N7139, N7140, N7141, N7049, N6587, OR4_1531_inw2, g38_inw1, N7624, N7489, N7626, N5145, N5069, N4515, N5059, N5058, N5310, N5071, N3834, N3988, N5309, N5073, N3835, N3989, N5239, N4267, N5308, N5075, N3836, N3990, N5307, N5077, N3837, N3991, N4978, N4979, N4976, N5057, N4027, N5162, N4199, N7703, AND4_1041_inw2, N3911, N5240, AND3_1508_inw1, AND3_1593_inw1, N3987, N5370, N5079, N3838, N3917, N5369, N5081, N3839, N3918, AND3_1022_inw1, AND3_1137_inw1, N4203, N5368, N5083, N3840, N3919, N5367, N5085, N3841, N3920, AND3_1138_inw1, N4200, N5311, N4523, N5366, N6835, N6837, N7871, N7873, N4357, OR4_1487_inw1, N4702, N4223, N5065, N6839, N6841, N7929, N7931, NOR3_1527_inw1, N4364, OR4_1526_inw1, N5364, N5106, N3908, N4701, N4224, N5363, N5108, N3909, N5140, N5110, N3914, N3975, N5371, N5305, N4521, N6162, N6160, AND4_1394_inw2, N5137, N6999, N7723, N7782, N4405, g16_inw1, N5304, N5115, N5303, N5113, N5306, N4855, N3915, N3976, AND3_840_inw1, AND3_1003_inw1, N4191, N3916, N3977, AND3_1004_inw1, N4188, NOR3_1524_invw, OR4_1522_inw2, N6100, N7080, N6896, N6097, N6138, AND3_1374_inw1, AND4_1368_inw1, N7787, N7788, N6651, n_305, N7076, N6890, N4733, AND3_1507_inw1, AND3_1590_inw1, N4524, NOR4_1525_invw, g30_inw2, g53_inw2, AND3_1340_inw1, N6099, AND4_1368_inw2, N6947, N8031, N8032, N6668, g2_inw1, g12_inw2, N4736, N5155, N4968, g10_inw1, N6504, N6536, AND3_1348_inw1, AND4_1341_inw1, AND4_1345_inw1, AND4_1349_inw2, N6948, N7984, N7985, N6670, g8_inw1, n_307, g32_inw1, N4735, N5154, N4965, N6096, N7218, N6897, N6891, N6133, N6949, N7851, N7852, N6672, g8_inw2, N4734, N5153, N4966, N6084, N6073, N6940, N7212, N6662, N7075, N6089, N7176, AND3_1332_inw1, AND4_1329_inw1, N7743, N7744, N6079, N6939, N7209, N6660, N7073, N4730, N5232, N5053, g10_inw2, N6946, N7917, N7918, N6666, g2_inw2, N4729, N5156, N4967, N6382, AND3_1321_inw1, AND4_1322_inw1, AND4_1329_inw2, N6935, N6936, N7879, N7880, N6653, N6066, N5241, NOR3_1513_invw, N6482, N6085, N6937, N6938, N7943, N7944, N6657, N4732, N6377, N5054, OR4_1486_inw2, N6814, N6411, N6490, N7815, N7816, N6661, N4731, N5233, N5052, OR4_1487_inw2, N7087, N6437, N6572, N6147, AND3_1383_inw1, AND4_1323_inw1, AND4_1381_inw2, N6689, N6691, N7821, N7822, N6690, N5235, N4725, N6143, N6074, N6958, N7222, N7181, AND4_1381_inw1, N7749, N7750, N6139, N6957, N7219, N7085, N5234, N4724, g14_inw2, AND3_1390_inw1, AND4_1391_inw1, N6964, N7887, N7923, N6695, g4_inw1, g6_inw2, N4728, N4975, N4974, NOR4_1538_invw, g26_inw2, g51_inw2, N6156, AND4_1414_inw2, N6965, N8009, N8034, N6434, n_303, g6_inw1, g16_inw2, N3827, g14_inw1, NOR3_1537_invw, N6584, N6606, AND3_1397_inw1, AND3_1419_inw1, AND4_1394_inw1, AND4_1398_inw2, AND4_1414_inw1, N6966, N7951, N7987, N6698, n_309, g28_inw1, N4727, N5161, N4972, N6154, N7229, N6916, N6909, N6194, N6189, N6699, N7823, N7859, N6700, g4_inw2, N4726, N5160, N4973, N8055, N8056, N8013, OR4_2241_inw1, OR4_1916_inw1, OR4_1974_inw1, OR4_1976_inw1, OR4_1977_inw1, OR4_1978_inw1, OR4_2088_inw1, OR4_2089_inw1, OR4_2090_inw1, OR4_2091_inw1, OR4_2300_inw1, N7505, N7727, N7728, N7729, N7730, N7435, N7507, N7508, N7509, N8121, OR4_1924_inw1, OR4_1979_inw1, OR4_1981_inw1, OR4_1982_inw1, OR4_1983_inw1, OR4_2092_inw1, OR4_2093_inw1, OR4_2094_inw1, OR4_2095_inw1, OR4_2301_inw1, N7510, N7731, N7732, N7733, N7734, N7443, N7512, N7513, N7514, N8122, N8057, N8058, N8017, OR4_2242_inw1, N4273, N4274, N4276, N4277, N7525, OR4_1992_inw1, N7449, N7736, N7737, N7738, N7739, N7515, N7516, N7517, N7518, N8123, OR4_1930_inw1, OR4_1987_inw1, OR4_1984_inw1, OR4_1985_inw1, OR4_1986_inw1, OR4_2097_inw1, OR4_2098_inw1, OR4_2099_inw1, OR4_2100_inw1, OR4_2302_inw1, OR4_1950_inw1, OR4_1988_inw1, OR4_1989_inw1, OR4_1990_inw1, OR4_1991_inw1, OR4_2096_inw1, OR4_2101_inw1, OR4_2102_inw1, OR4_2103_inw1, OR4_2303_inw1, N7735, N7740, N7741, N7742, N7519, N7520, N7521, N7522, N8124, N7469, N8075, N8076, OR3_1670_inw1, OR3_1837_inw1, OR3_1840_inw1, OR3_1867_inw1, OR3_1868_inw1, OR3_1869_inw1, OR3_1870_inw1, OR3_1871_inw1, OR3_1874_inw1, OR3_1875_inw1, OR3_1998_inw1, OR3_1999_inw1, OR3_2000_inw1, OR3_2001_inw1, OR3_2002_inw1, OR3_2003_inw1, OR3_2004_inw1, OR3_2005_inw1, OR4_2278_inw1, OR4_2279_inw1, N7365, N7473, N7472, N7471, N7015, N7363, N7467, N7466, N7470, N7707, N7706, N7705, N7704, N7465, N7702, N7701, N7700, N7699, N7037, N7245, N7236, N7239, N7242, N7173, N7174, N7175, N6828, N6827, g33_invw, N4278, N6967, N7263, N7250, N7257, N7260, N7178, N7179, N7180, N6855, N6854, g38_invw, N7698, N7625, N5711, N5385, N5707, N5703, N5331, N5332, N5163, N5164, N5236, N4721, N5328, N5060, N6475, N6722, AND3_1509_inw1, AND3_1592_inw1, N5742, AND3_1023_inw1, N5745, N5736, N7044, N7045, N7900, N7903, AND3_1046_inw1, N6953, N6954, N7885, N7886, N6386, N5049, N5365, N7046, N7047, N7960, N7963, NOR3_1527_invw, N6144, N6955, N6956, N7945, N7946, N6566, N5739, N5700, N6024, N6023, N5696, OR4_1535_inw2, N6157, N7090, N7778, N7812, N6915, N7751, N7795, N6155, N5692, AND3_1005_inw1, N6553, NOR4_1525_inw2, g30_inw1, g53_inw1, N7217, N6127, N7800, N7803, N7769, N7771, N7216, N7215, AND4_1044_inw1, N6474, N6719, AND3_1506_inw1, AND3_1591_inw1, N6556, N6500, N6539, N7031, N8037, N8038, N6826, N8021, N8023, N6117, AND4_1044_inw2, N5319, N6397, N6825, N6889, N7034, N7998, N8001, N7967, N7969, N6091, N5315, N7412, N7321, N7320, N7079, N7864, N7867, N7833, N7835, OR4_1512_inw2, N7408, N7407, N6881, N6080, N7762, N7765, N7709, N7711, N7022, N7406, N7405, AND4_1043_inw1, N5377, N7028, N7932, N7935, N6824, N7897, N7899, N6924, N7018, N7019, N7890, N7893, N6808, N6810, N7861, N7863, N6634, N5388, N6486, N7492, N6807, N7020, N7021, N7954, N7957, N6812, N7925, N7927, AND4_1043_inw2, N6811, N7826, N7829, N7797, N7799, N6901, N6838, N6140, N7836, N7839, N7807, N7809, N5382, AND4_1041_inw1, OR4_1526_inw2, N7418, N7417, N7772, N7775, N7719, N7721, N7048, N7416, N7415, N6427, N7054, N7906, N7940, N6851, N7875, N7910, N6149, N6175, AND4_1042_inw2, N6622, N6580, N6609, NOR4_1538_inw2, g26_inw1, g51_inw1, N6184, N7057, N8025, N8039, N6853, N7993, N8027, N6619, N6852, N7160, N6912, N7060, N7970, N8004, N7939, N7974, AND4_1042_inw1, N5324, N7421, N7328, N7089, N7088, N7842, N7876, N7811, N7846, N8061, N8059, N8033, N8064, N8060, N8036, n_320, n_321, n_318, n_325, N7432, n_322, n_323, N6714, N6715, N6710, N6477, N6044, AND3_1586_inw1, AND3_1668_inw1, N6206, AND3_1669_inw1, N6203, N5756, N6378, N5755, N6476, N6471, AND3_1175_inw1, N6874, N6875, N6721, N6633, N6375, N6632, N6376, N6631, N6373, N7130, N7928, N7930, N6925, N6221, N5312, N7131, AND3_2234_inw1, AND3_2236_inw1, AND3_2233_inw1, AND3_2235_inw1, N6569, N7498, N6834, N6630, N6374, N6712, N6713, N6708, N6716, AND3_1584_inw1, AND3_1666_inw1, N6200, N7228, N7810, N7845, AND3_1667_inw1, N6197, N6895, N7832, N7834, N7409, N5063, N6873, N6872, N6473, N6720, N7658, N6900, N6823, N7657, N6894, n_319, N8040, N6641, N6675, N6469, N6801, AND3_2228_inw1, N6831, N8020, N8022, N6648, N6025, N7588, N7587, N7896, N7898, N7582, N7493, N7072, N7796, N7798, N7579, N5062, N7002, N6067, N7966, N7968, N6926, N7115, N7924, N7926, N6923, N6922, N6809, N7116, AND3_2230_inw1, AND3_2227_inw1, AND3_2229_inw1, N7860, N7862, N7084, N6643, N6646, N6802, N7870, N7872, N6069, N6068, N7592, N7499, N7806, N7808, N7589, N6857, n_324, N7938, N7973, N6703, N5061, N7665, N6919, N6850, N7500, N6913, N8042, N6914, N7225, N7992, N8026, N6028, N7599, N7598, N7874, N7909, N8073, N8074, g37_inw2, g37_inw1, g43_inw2, n_326, g43_inw1, N6975, N6976, N6862, N6863, N6877, N6235, AND3_1587_inw1, N6234, N6637, N7006, N6795, N6792, N6927, N6836, N6973, N6974, N6860, N6861, g44_invw, AND3_1585_inw1, N7586, N7585, AND3_1237_inw1, N7003, N7715, N7712, N7041, N7710, N7708, N7101, N7720, N7718, N7065, N7724, N7595, N7420, N7419, N7503, N7504, N7097, n_327, N7206, N6876, N7151, N7150, N7269, N6978, N7268, N6977, N7094, n_328, N7300, N7149, N7770, N7768, N7177, N7204, N7205, N7182, N7781, N7722, N7186, N7185, N7301, N7476, N7474, N7184, N7183, N7402, N7468, g44_inw1, N7529;
	wire g44_inw1_key, N7402_key, N7184_key, N7474_key, N7476_key, N7301_key, N7186_key, N7204_key, N7300_key, N7094_key, N7268_key, N7269_key, N372_key, N2954_key, N3723_key, N4008_key, N5366_key, N5364_key, N5363_key, N5140_key, N5305_key, N5137_key, N5304_key, N5303_key, N5306_key, N5736_key, N5739_key, N5700_key, N5696_key, N5692_key, N6631_key, N6630_key, N6712_key, N6713_key, AND3_1584_inw1_key, AND3_1666_inw1_key, AND3_1667_inw1_key, N6792_key, N6973_key, N6974_key, N6860_key, N6861_key, AND3_1585_inw1_key, N292_key, N3680_key, N2867_key, N4011_key, N5145_key, N5310_key, N5309_key, N5308_key, N5307_key, N5370_key, N5369_key, N5368_key, N5367_key, N5311_key, N5711_key, N5707_key, N5703_key, N5742_key, N5745_key, N6714_key, N6715_key, AND3_1586_inw1_key, AND3_1668_inw1_key, AND3_1669_inw1_key, N6633_key, N6632_key, N6975_key, N6976_key, N6862_key, N6863_key, AND3_1587_inw1_key, N6795_key, N7097_key, N566_key, N3027_key, N3023_key, N3028_key, N3024_key, N3029_key, N3025_key, N3030_key, N3026_key, N2938_key, N2939_key, N2940_key, N2941_key, AND3_377_inw1_key, AND3_378_inw1_key, AND3_379_inw1_key, AND3_380_inw1_key, AND3_444_inw1_key, AND3_445_inw1_key, AND3_446_inw1_key, AND3_447_inw1_key, AND3_524_inw1_key, AND3_525_inw1_key, AND3_526_inw1_key, AND3_527_inw1_key, AND3_547_inw1_key, AND3_548_inw1_key, AND3_549_inw1_key, AND3_550_inw1_key, N3463_key, N3464_key, N3465_key, N3466_key, N3508_key, N3509_key, N3510_key, N3511_key, N2934_key, N2935_key, N2936_key, N2937_key, N4608_key, N3722_key, N3719_key, N3720_key, N3721_key, N3769_key, N3770_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123;
	assign N3360 = N1;
	assign N3359 = N1;
	assign N3358 = N1;
	assign N3357 = N1;
	assign N2309 = N1;
	assign N1146 = ~( N373 & N1 );
	assign N6107 = ( N4 & N5462 );
	assign N6664 = ( N6091 & N4 );
	assign AND3_1351_inw1 = ~( N4 & N5462 );
	assign AND4_1349_inw1 = ~( N4 & N5462 );
	assign N6806 = ~( N4 & N6651 );
	assign N2637 = ~N4;
	assign AND3_600_inw1 = ~( N11 & N2779 );
	assign AND3_619_inw1 = ~( N11 & N2801 );
	assign AND3_609_inw1 = ~( N14 & N2779 );
	assign AND3_617_inw1 = ~( N14 & N2801 );
	assign AND3_230_inw1 = ~( N17 & N610 );
	assign AND3_238_inw1 = ~( N17 & N613 );
	assign AND3_229_inw1 = ~( N20 & N610 );
	assign AND3_237_inw1 = ~( N20 & N613 );
	assign AND3_813_inw1 = ~( N23 & N588 );
	assign AND3_807_inw1 = ~( N24 & N1588 );
	assign AND3_808_inw1 = ~( N25 & N588 );
	assign AND3_809_inw1 = ~( N26 & N1588 );
	assign N1150 = ( N1043 & N27 );
	assign N1475 = ( N27 & N31 );
	assign N3740 = ( N34 & N588 );
	assign AND3_228_inw1 = ~( N37 & N610 );
	assign AND3_236_inw1 = ~( N37 & N613 );
	assign AND3_227_inw1 = ~( N40 & N610 );
	assign AND3_235_inw1 = ~( N40 & N613 );
	assign AND3_605_inw1 = ~( N43 & N2779 );
	assign AND3_613_inw1 = ~( N43 & N2801 );
	assign AND3_602_inw1 = ~( N46 & N2779 );
	assign AND3_610_inw1 = ~( N46 & N2801 );
	assign AND3_225_inw1 = ~( N49 & N610 );
	assign AND3_233_inw1 = ~( N49 & N613 );
	assign AND3_733_inw1 = ~( N52 & N3068 );
	assign AND3_730_inw1 = ~( N53 & N3068 );
	assign N5119 = ( N54 & N4405 );
	assign N6693 = ( N6149 & N54 );
	assign AND3_1400_inw1 = ~( N54 & N4405 );
	assign AND4_1398_inw1 = ~( N54 & N4405 );
	assign N5955 = ~( N54 & N3921 );
	assign N2715 = ~N54;
	assign AND3_223_inw1 = ~( N61 & N610 );
	assign AND3_244_inw1 = ~( N61 & N613 );
	assign AND3_232_inw1 = ~( N64 & N610 );
	assign AND3_240_inw1 = ~( N64 & N613 );
	assign AND3_608_inw1 = ~( N67 & N2779 );
	assign AND3_616_inw1 = ~( N67 & N2801 );
	assign AND3_231_inw1 = ~( N70 & N610 );
	assign AND3_239_inw1 = ~( N70 & N613 );
	assign AND3_607_inw1 = ~( N73 & N2779 );
	assign AND3_615_inw1 = ~( N73 & N2801 );
	assign AND3_606_inw1 = ~( N76 & N2779 );
	assign AND3_614_inw1 = ~( N76 & N2801 );
	assign AND3_812_inw1 = ~( N79 & N1588 );
	assign AND3_815_inw1 = ~( N80 & N588 );
	assign AND3_810_inw1 = ~( N81 & N588 );
	assign AND3_814_inw1 = ~( N82 & N1588 );
	assign N2969 = ( N83 & N1588 );
	assign N3738 = ( N83 & N588 );
	assign N2970 = ( N86 & N1588 );
	assign N3739 = ( N87 & N588 );
	assign N2971 = ( N88 & N1588 );
	assign AND3_604_inw1 = ~( N91 & N2779 );
	assign AND3_612_inw1 = ~( N91 & N2801 );
	assign N3072 = ( N94 & N625 );
	assign N3071 = ( N97 & N625 );
	assign AND3_603_inw1 = ~( N100 & N2779 );
	assign AND3_611_inw1 = ~( N100 & N2801 );
	assign AND3_226_inw1 = ~( N103 & N610 );
	assign AND3_234_inw1 = ~( N103 & N613 );
	assign AND3_222_inw1 = ~( N106 & N613 );
	assign AND3_224_inw1 = ~( N106 & N610 );
	assign AND3_597_inw1 = ~( N109 & N2801 );
	assign AND3_601_inw1 = ~( N109 & N2779 );
	assign AND3_734_inw1 = ~( N112 & N3068 );
	assign AND3_729_inw1 = ~( N113 & N3068 );
	assign AND3_731_inw1 = ~( N114 & N3068 );
	assign AND3_732_inw1 = ~( N115 & N3068 );
	assign AND3_735_inw1 = ~( N116 & N3068 );
	assign AND3_717_inw1 = ~( N117 & N3068 );
	assign AND3_620_inw1 = ~( N118 & N3068 );
	assign AND3_723_inw1 = ~( N119 & N3068 );
	assign AND3_618_inw1 = ~( N120 & N3068 );
	assign AND3_736_inw1 = ~( N121 & N3068 );
	assign AND3_728_inw1 = ~( N122 & N3068 );
	assign AND3_242_inw1 = ~( N123 & N1758 );
	assign AND3_737_inw1 = ~( N123 & N3068 );
	assign AND3_718_inw1 = ~( N126 & N3068 );
	assign AND3_719_inw1 = ~( N127 & N3068 );
	assign AND3_720_inw1 = ~( N128 & N3068 );
	assign AND3_722_inw1 = ~( N129 & N3068 );
	assign AND3_724_inw1 = ~( N130 & N3068 );
	assign AND3_721_inw1 = ~( N131 & N3068 );
	assign N6880 = ( N6478 & N132 );
	assign N6478 = ~( N4357 & N132 );
	assign N1042 = ( N135 & N631 );
	assign N2054 = ( N136 & N1148 );
	assign N2139 = N137;
	assign N7506 = ( N7435 & N137 );
	assign N7511 = ( N7443 & N137 );
	assign N7600 = ( N7505 & N137 );
	assign N7601 = ( N7507 & N137 );
	assign N7602 = ( N7508 & N137 );
	assign N7603 = ( N7509 & N137 );
	assign N7604 = ( N7510 & N137 );
	assign N7605 = ( N7512 & N137 );
	assign N7606 = ( N7513 & N137 );
	assign N7607 = ( N7514 & N137 );
	assign N7754 = ( N7727 & N137 );
	assign N7755 = ( N7728 & N137 );
	assign N7756 = ( N7729 & N137 );
	assign N7757 = ( N7730 & N137 );
	assign N7758 = ( N7731 & N137 );
	assign N7759 = ( N7732 & N137 );
	assign N7760 = ( N7733 & N137 );
	assign N7761 = ( N7734 & N137 );
	assign N8125 = ( N8121 & N137 );
	assign N8126 = ( N8122 & N137 );
	assign N2590 = ~( N1475 & N140 );
	assign N2142 = N141;
	assign N709 = N141;
	assign N1147 = ( N141 & N145 );
	assign N4737 = ( N4273 & N141 );
	assign N4738 = ( N4274 & N141 );
	assign N4739 = ( N4276 & N141 );
	assign N4740 = ( N4277 & N141 );
	assign AND3_212_inw1 = ~( N146 & N571 );
	assign AND3_221_inw1 = ~( N146 & N577 );
	assign AND3_583_inw1 = ~( N149 & N2653 );
	assign AND3_594_inw1 = ~( N149 & N2728 );
	assign AND3_211_inw1 = ~( N152 & N571 );
	assign AND3_220_inw1 = ~( N152 & N577 );
	assign AND3_582_inw1 = ~( N155 & N2653 );
	assign AND3_593_inw1 = ~( N155 & N2728 );
	assign AND3_210_inw1 = ~( N158 & N571 );
	assign AND3_219_inw1 = ~( N158 & N577 );
	assign AND3_207_inw1 = ~( N161 & N571 );
	assign AND3_217_inw1 = ~( N161 & N577 );
	assign AND3_206_inw1 = ~( N164 & N571 );
	assign AND3_216_inw1 = ~( N164 & N577 );
	assign AND3_205_inw1 = ~( N167 & N571 );
	assign AND3_215_inw1 = ~( N167 & N577 );
	assign AND3_203_inw1 = ~( N170 & N571 );
	assign AND3_213_inw1 = ~( N170 & N577 );
	assign AND3_204_inw1 = ~( N173 & N571 );
	assign AND3_214_inw1 = ~( N173 & N577 );
	assign AND3_621_inw1 = ~( N176 & N2653 );
	assign AND3_622_inw1 = ~( N176 & N2728 );
	assign AND3_271_inw1 = ~( N179 & N571 );
	assign AND3_292_inw1 = ~( N179 & N577 );
	assign AND3_580_inw1 = ~( N182 & N2653 );
	assign AND3_591_inw1 = ~( N182 & N2728 );
	assign AND3_209_inw1 = ~( N185 & N571 );
	assign AND3_218_inw1 = ~( N185 & N577 );
	assign AND3_581_inw1 = ~( N188 & N2653 );
	assign AND3_592_inw1 = ~( N188 & N2728 );
	assign AND3_579_inw1 = ~( N191 & N2653 );
	assign AND3_590_inw1 = ~( N191 & N2728 );
	assign AND3_578_inw1 = ~( N194 & N2653 );
	assign AND3_589_inw1 = ~( N194 & N2728 );
	assign AND3_577_inw1 = ~( N197 & N2653 );
	assign AND3_588_inw1 = ~( N197 & N2728 );
	assign AND3_575_inw1 = ~( N200 & N2653 );
	assign AND3_586_inw1 = ~( N200 & N2728 );
	assign AND3_576_inw1 = ~( N203 & N2653 );
	assign AND3_587_inw1 = ~( N203 & N2728 );
	assign N3689 = ( N206 & N2855 );
	assign N3761 = ( N242 & N206 );
	assign N3758 = ~( AND3_700_inw1 | N206 );
	assign N3823 = ~( N206 & N2823 );
	assign N3753 = ~N206;
	assign N2876 = ( N209 & N335 );
	assign N2835 = ( N1067 & N210 );
	assign N3027 = ( N242 & N210 );
	assign N3688 = ( N210 & N2855 );
	assign N2831 = ~( AND3_305_inw1 | N210 );
	assign N3023 = ~( AND3_444_inw1_key | N210 );
	assign N4024 = ~( N210 & N3753 );
	assign N2823 = ~N210;
	assign N2875 = ( N217 & N335 );
	assign N2836 = ( N1067 & N218 );
	assign N3028 = ( N242 & N218 );
	assign N3687 = ( N218 & N2855 );
	assign N2832 = ~( AND3_306_inw1 | N218 );
	assign N3024 = ~( AND3_445_inw1_key | N218 );
	assign N3610 = ~( N218 & N2827 );
	assign N2825 = ~N218;
	assign N2874 = ( N225 & N335 );
	assign N2837 = ( N1067 & N226 );
	assign N3029 = ( N242 & N226 );
	assign N3686 = ( N226 & N2855 );
	assign N2833 = ~( AND3_307_inw1 | N226 );
	assign N3025 = ~( AND3_446_inw1_key | N226 );
	assign N3609 = ~( N226 & N2825 );
	assign N2827 = ~N226;
	assign N2873 = ( N233 & N335 );
	assign N2838 = ( N1067 & N234 );
	assign N3030 = ( N242 & N234 );
	assign N3685 = ( N234 & N2855 );
	assign N2834 = ~( AND3_308_inw1 | N234 );
	assign N3026 = ~( AND3_447_inw1_key | N234 );
	assign N3563 = ~( N234 & N2839 );
	assign N2829 = ~N234;
	assign N2872 = ( N241 & N335 );
	assign N2910 = ( N242 & N293 );
	assign N2911 = ( N242 & N308 );
	assign N2912 = ( N242 & N316 );
	assign N2938 = ( N242 & N257 );
	assign N2939 = ( N242 & N265 );
	assign N2940 = ( N242 & N273 );
	assign N2941 = ( N242 & N281 );
	assign N2983 = ( N242 & N324 );
	assign N2985 = ( N242 & N341 );
	assign N2986 = ( N242 & N351 );
	assign N2984 = ( N242 | N514 );
	assign N1152 = ~N245;
	assign n_331 = ( N562 & N245 );
	assign N2907 = ( N248 & N302 );
	assign N2980 = ( N248 & N514 );
	assign N3013 = ( N248 & N361 );
	assign AND3_351_inw1 = ~( N248 & N479 );
	assign AND3_352_inw1 = ~( N248 & N490 );
	assign AND3_377_inw1 = ~( N248 & N389 );
	assign AND3_378_inw1 = ~( N248 & N400 );
	assign AND3_379_inw1 = ~( N248 & N411 );
	assign AND3_380_inw1 = ~( N248 & N374 );
	assign AND3_408_inw1 = ~( N248 & N503 );
	assign AND3_410_inw1 = ~( N248 & N523 );
	assign AND3_411_inw1 = ~( N248 & N534 );
	assign AND3_444_inw1 = ~( N248 & N457 );
	assign AND3_445_inw1 = ~( N248 & N468 );
	assign AND3_446_inw1 = ~( N248 & N422 );
	assign AND3_447_inw1 = ~( N248 & N435 );
	assign AND3_700_inw1 = ~( N248 & N446 );
	assign N3444 = ( N251 & N2902 );
	assign N3502 = ( N251 & N2999 );
	assign AND3_512_inw1 = ~( N479 & N251 );
	assign AND3_513_inw1 = ~( N490 & N251 );
	assign AND3_524_inw1 = ~( N389 & N251 );
	assign AND3_525_inw1 = ~( N400 & N251 );
	assign AND3_526_inw1 = ~( N411 & N251 );
	assign AND3_527_inw1 = ~( N374 & N251 );
	assign AND3_532_inw1 = ~( N503 & N251 );
	assign AND3_534_inw1 = ~( N523 & N251 );
	assign AND3_535_inw1 = ~( N534 & N251 );
	assign AND3_547_inw1 = ~( N457 & N251 );
	assign AND3_548_inw1 = ~( N468 & N251 );
	assign AND3_549_inw1 = ~( N422 & N251 );
	assign AND3_550_inw1 = ~( N435 & N251 );
	assign AND3_790_inw1 = ~( N446 & N251 );
	assign N3447 = ( N254 & N2901 );
	assign N3448 = ( N254 & N2903 );
	assign N3449 = ( N254 & N2905 );
	assign N3463 = ( N254 & N2839 );
	assign N3464 = ( N254 & N2841 );
	assign N3465 = ( N254 & N2843 );
	assign N3466 = ( N254 & N2845 );
	assign N3485 = ( N254 & N1660 );
	assign N3486 = ( N254 & N2915 );
	assign N3487 = ( N254 & N2917 );
	assign N3508 = ( N254 & N2823 );
	assign N3509 = ( N254 & N2825 );
	assign N3510 = ( N254 & N2827 );
	assign N3511 = ( N254 & N2829 );
	assign N3982 = ( N254 & N3753 );
	assign N2851 = ( N1067 & N257 );
	assign N3684 = ( N257 & N2855 );
	assign N2847 = ~( AND3_321_inw1 | N257 );
	assign N2934 = ~( AND3_377_inw1_key | N257 );
	assign N3562 = ~( N257 & N2829 );
	assign N2839 = ~N257;
	assign N2871 = ( N264 & N335 );
	assign N2852 = ( N1067 & N265 );
	assign N3683 = ( N265 & N2855 );
	assign N2848 = ~( AND3_322_inw1 | N265 );
	assign N2935 = ~( AND3_378_inw1_key | N265 );
	assign N3561 = ~( N265 & N2843 );
	assign N2841 = ~N265;
	assign N2870 = ( N272 & N335 );
	assign N2853 = ( N1067 & N273 );
	assign N3682 = ( N273 & N2855 );
	assign N2849 = ~( AND3_323_inw1 | N273 );
	assign N2936 = ~( AND3_379_inw1_key | N273 );
	assign N3560 = ~( N273 & N2841 );
	assign N2843 = ~N273;
	assign N2869 = ( N280 & N335 );
	assign N2854 = ( N1067 & N281 );
	assign N3681 = ( N281 & N2855 );
	assign N2850 = ~( AND3_324_inw1 | N281 );
	assign N2937 = ~( AND3_380_inw1_key | N281 );
	assign N3559 = ~( N281 & N3142 );
	assign N2845 = ~N281;
	assign N2868 = ( N288 & N335 );
	assign N3680 = ( N289 & N2855 );
	assign N3558 = ~( N289 & N2845 );
	assign N3142 = ~N289;
	assign N2867 = ( N292_key & N335 );
	assign N816 = N293;
	assign N3731 = ( N293 & N2942 );
	assign N3608 = ~( N293 & N2902 );
	assign N2901 = ~N293;
	assign N3604 = N299;
	assign N2527 = N299;
	assign N2963 = ( N299 & N332 );
	assign N3613 = ~N299;
	assign N3730 = ( N302 & N2942 );
	assign N3607 = ~( N302 & N2901 );
	assign N2902 = ~N302;
	assign N2962 = ( N307 & N332 );
	assign N3729 = ( N308 & N2942 );
	assign N2908 = ~( AND3_351_inw1 | N308 );
	assign N3606 = ~( N308 & N2905 );
	assign N2903 = ~N308;
	assign N2961 = ( N315 & N332 );
	assign N3728 = ( N316 & N2942 );
	assign N2909 = ~( AND3_352_inw1 | N316 );
	assign N3605 = ~( N316 & N2903 );
	assign N2905 = ~N316;
	assign N2960 = ( N323 & N332 );
	assign N2923 = ( N1067 & N324 );
	assign N3727 = ( N324 & N2942 );
	assign N2919 = ~( AND3_362_inw1 | N324 );
	assign N2979 = ~( AND3_408_inw1 | N324 );
	assign N4953 = ~( AND3_1003_inw1 | N324 );
	assign N4954 = ~( AND3_1004_inw1 | N324 );
	assign N1660 = ~N324;
	assign N2959 = ( N331 & N332 );
	assign N2954 = ( N372_key & N332 );
	assign N2955 = ( N366 & N332 );
	assign N2956 = ( N358 & N332 );
	assign N2957 = ( N348 & N332 );
	assign N2958 = ( N338 & N332 );
	assign N2942 = ~N332;
	assign N2855 = ~N335;
	assign N1144 = ~N338;
	assign N2924 = ( N1067 & N341 );
	assign N3726 = ( N341 & N2942 );
	assign N2921 = ~( AND3_364_inw1 | N341 );
	assign N2981 = ~( AND3_410_inw1 | N341 );
	assign N3515 = ~( N341 & N2917 );
	assign N2915 = ~N341;
	assign N1138 = ~N348;
	assign N2925 = ( N1067 & N351 );
	assign N3725 = ( N351 & N2942 );
	assign N2922 = ~( AND3_365_inw1 | N351 );
	assign N2982 = ~( AND3_411_inw1 | N351 );
	assign N3514 = ~( N351 & N2915 );
	assign N2917 = ~N351;
	assign N1145 = ~N358;
	assign N3724 = ( N361 & N2942 );
	assign N3513 = ~( N361 & N3032 );
	assign N2999 = ~N361;
	assign N1139 = ~N366;
	assign N3723 = ( N369 & N2942 );
	assign N3512 = ~( N369 & N2999 );
	assign N3032 = ~N369;
	assign N4310 = ( N3842 & N374 );
	assign AND3_324_inw1 = ~( N1104 & N374 );
	assign AND3_506_inw1 = ~( N374 & N1092 );
	assign N5250 = ~( N374 & N5085 );
	assign N4608 = ~( N374 | N3842 );
	assign N2636 = ~N374;
	assign N3679 = ~( OR3_638_inw1 & N374 );
	assign N3722 = ~( OR3_669_inw1 & N374 );
	assign N1151 = ( N386 & N556 );
	assign g45_inw1 = ~( n_327 & N386 );
	assign N4298 = ( N3861 & N389 );
	assign AND3_321_inw1 = ~( N1104 & N389 );
	assign AND3_503_inw1 = ~( N389 & N1092 );
	assign N5247 = ~( N389 & N5079 );
	assign N2633 = ~N389;
	assign N3676 = ~( OR3_635_inw1 & N389 );
	assign N3719 = ~( OR3_666_inw1 & N389 );
	assign N4301 = ( N3855 & N400 );
	assign AND3_322_inw1 = ~( N1104 & N400 );
	assign AND3_504_inw1 = ~( N400 & N1092 );
	assign N5248 = ~( N400 & N5081 );
	assign N2634 = ~N400;
	assign N3677 = ~( OR3_636_inw1 & N400 );
	assign N3720 = ~( OR3_667_inw1 & N400 );
	assign N4305 = ( N3849 & N411 );
	assign AND3_323_inw1 = ~( N1104 & N411 );
	assign AND3_505_inw1 = ~( N411 & N1092 );
	assign N5249 = ~( N411 & N5083 );
	assign N2635 = ~N411;
	assign N3678 = ~( OR3_637_inw1 & N411 );
	assign N3721 = ~( OR3_668_inw1 & N411 );
	assign N4290 = ( N422 & N3873 );
	assign AND3_307_inw1 = ~( N1104 & N422 );
	assign AND3_497_inw1 = ~( N422 & N1092 );
	assign N5245 = ~( N422 & N5075 );
	assign N4575 = ~( N422 | N3873 );
	assign N2631 = ~N422;
	assign N3670 = ~( OR3_629_inw1 & N422 );
	assign N3769 = ~( OR3_711_inw1 & N422 );
	assign N4297 = ( N3867 & N435 );
	assign AND3_308_inw1 = ~( N1104 & N435 );
	assign AND3_498_inw1 = ~( N435 & N1092 );
	assign N5246 = ~( N435 & N5077 );
	assign N2632 = ~N435;
	assign N3671 = ~( OR3_630_inw1 & N435 );
	assign N3770 = ~( OR3_712_inw1 & N435 );
	assign N4268 = ( N446 & N3893 );
	assign N5242 = ~( N446 & N5069 );
	assign N2628 = ~N446;
	assign N4185 = ~( OR3_836_inw1 & N446 );
	assign N4280 = ( N3887 & N457 );
	assign AND3_305_inw1 = ~( N1104 & N457 );
	assign AND3_495_inw1 = ~( N457 & N1092 );
	assign N5243 = ~( N457 & N5071 );
	assign N2629 = ~N457;
	assign N3668 = ~( OR3_627_inw1 & N457 );
	assign N3767 = ~( OR3_709_inw1 & N457 );
	assign N4284 = ( N3881 & N468 );
	assign AND3_306_inw1 = ~( N1104 & N468 );
	assign AND3_496_inw1 = ~( N468 & N1092 );
	assign N5244 = ~( N468 & N5073 );
	assign N2630 = ~N468;
	assign N3669 = ~( OR3_628_inw1 & N468 );
	assign N3768 = ~( OR3_710_inw1 & N468 );
	assign N4379 = ( N3956 & N479 );
	assign N5261 = ~( N479 & N5106 );
	assign N2709 = ~N479;
	assign N3703 = ~( OR3_653_inw1 & N479 );
	assign N4385 = ( N490 & N3948 );
	assign N5262 = ~( N490 & N5108 );
	assign N4627 = ~( N490 | N3948 );
	assign N2710 = ~N490;
	assign N3704 = ~( OR3_654_inw1 & N490 );
	assign N4392 = ( N3942 & N503 );
	assign AND3_362_inw1 = ~( N1104 & N503 );
	assign AND3_517_inw1 = ~( N503 & N1092 );
	assign N5263 = ~( N503 & N5110 );
	assign N2711 = ~N503;
	assign N3711 = ~( OR3_659_inw1 & N503 );
	assign N3745 = ~( OR3_687_inw1 & N503 );
	assign N2349 = ( N1104 & N514 );
	assign N4067 = ( N3732 & N514 );
	assign N5112 = ~( N514 & N4855 );
	assign N2712 = ~N514;
	assign N2350 = ( N1067 | N514 );
	assign N4396 = ( N3933 & N523 );
	assign AND3_364_inw1 = ~( N1104 & N523 );
	assign AND3_518_inw1 = ~( N523 & N1092 );
	assign N5274 = ~( N523 & N5113 );
	assign N2713 = ~N523;
	assign N3712 = ~( OR3_660_inw1 & N523 );
	assign N3746 = ~( OR3_688_inw1 & N523 );
	assign N4400 = ( N3927 & N534 );
	assign AND3_365_inw1 = ~( N1104 & N534 );
	assign AND3_519_inw1 = ~( N534 & N1092 );
	assign N5275 = ~( N534 & N5115 );
	assign N2714 = ~N534;
	assign N3713 = ~( OR3_661_inw1 & N534 );
	assign N3747 = ~( OR3_689_inw1 & N534 );
	assign N1137 = ~N545;
	assign N2387 = N549;
	assign N1141 = ~N549;
	assign N1140 = ( N552 & N562 );
	assign N1153 = ~N552;
	assign n_330 = ( N556 & N552 );
	assign N1155 = ~N559;
	assign n_329 = ~( g45_inw1 | N559 );
	assign N1154 = ~N562;
	assign N8041 = ( N566_key & N8037 );
	assign N7990 = ~( AND3_2229_inw1 | N566_key );
	assign N7991 = ~( AND3_2230_inw1 | N566_key );
	assign N1157 = ~N566_key;
	assign AND3_1879_inw1 = ~( N7190 & N571 );
	assign AND3_1915_inw1 = ~( N7304 & N571 );
	assign AND3_1917_inw1 = ~( N7270 & N571 );
	assign AND3_1919_inw1 = ~( N7276 & N571 );
	assign AND3_1921_inw1 = ~( N7282 & N571 );
	assign AND3_2034_inw1 = ~( N7531 & N571 );
	assign AND3_2036_inw1 = ~( N7537 & N571 );
	assign AND3_2038_inw1 = ~( N7543 & N571 );
	assign AND3_2040_inw1 = ~( N7549 & N571 );
	assign AND3_2297_inw1 = ~( N8093 & N571 );
	assign N2653 = ~N571;
	assign N2585 = ~( AND3_203_inw1 | N574 );
	assign N2586 = ~( AND3_204_inw1 | N574 );
	assign N2587 = ~( AND3_205_inw1 | N574 );
	assign N2588 = ~( AND3_206_inw1 | N574 );
	assign N2589 = ~( AND3_207_inw1 | N574 );
	assign N2591 = ~( AND3_209_inw1 | N574 );
	assign N2592 = ~( AND3_210_inw1 | N574 );
	assign N2593 = ~( AND3_211_inw1 | N574 );
	assign N2594 = ~( AND3_212_inw1 | N574 );
	assign N2703 = ~( AND3_271_inw1 | N574 );
	assign N3616 = ~( AND3_575_inw1 | N574 );
	assign N3617 = ~( AND3_576_inw1 | N574 );
	assign N3618 = ~( AND3_577_inw1 | N574 );
	assign N3619 = ~( AND3_578_inw1 | N574 );
	assign N3620 = ~( AND3_579_inw1 | N574 );
	assign N3621 = ~( AND3_580_inw1 | N574 );
	assign N3622 = ~( AND3_581_inw1 | N574 );
	assign N3623 = ~( AND3_582_inw1 | N574 );
	assign N3624 = ~( AND3_583_inw1 | N574 );
	assign N3662 = ~( AND3_621_inw1 | N574 );
	assign N2664 = ~N574;
	assign AND3_1881_inw1 = ~( N7190 & N577 );
	assign AND3_1923_inw1 = ~( N7304 & N577 );
	assign AND3_1925_inw1 = ~( N7270 & N577 );
	assign AND3_1927_inw1 = ~( N7276 & N577 );
	assign AND3_1929_inw1 = ~( N7282 & N577 );
	assign AND3_2042_inw1 = ~( N7531 & N577 );
	assign AND3_2044_inw1 = ~( N7537 & N577 );
	assign AND3_2046_inw1 = ~( N7543 & N577 );
	assign AND3_2048_inw1 = ~( N7549 & N577 );
	assign AND3_2299_inw1 = ~( N8093 & N577 );
	assign N2728 = ~N577;
	assign N2595 = ~( AND3_213_inw1 | N580 );
	assign N2596 = ~( AND3_214_inw1 | N580 );
	assign N2597 = ~( AND3_215_inw1 | N580 );
	assign N2598 = ~( AND3_216_inw1 | N580 );
	assign N2599 = ~( AND3_217_inw1 | N580 );
	assign N2600 = ~( AND3_218_inw1 | N580 );
	assign N2601 = ~( AND3_219_inw1 | N580 );
	assign N2602 = ~( AND3_220_inw1 | N580 );
	assign N2603 = ~( AND3_221_inw1 | N580 );
	assign N2778 = ~( AND3_292_inw1 | N580 );
	assign N3627 = ~( AND3_586_inw1 | N580 );
	assign N3628 = ~( AND3_587_inw1 | N580 );
	assign N3629 = ~( AND3_588_inw1 | N580 );
	assign N3630 = ~( AND3_589_inw1 | N580 );
	assign N3631 = ~( AND3_590_inw1 | N580 );
	assign N3632 = ~( AND3_591_inw1 | N580 );
	assign N3633 = ~( AND3_592_inw1 | N580 );
	assign N3634 = ~( AND3_593_inw1 | N580 );
	assign N3635 = ~( AND3_594_inw1 | N580 );
	assign N3663 = ~( AND3_622_inw1 | N580 );
	assign N2739 = ~N580;
	assign N8035 = ( N583 & N8025 );
	assign N7996 = ~( AND3_2235_inw1 | N583 );
	assign N7997 = ~( AND3_2236_inw1 | N583 );
	assign N1219 = ~N583;
	assign N3615 = ( N588 & N2623 );
	assign N1588 = ~N588;
	assign N1043 = ~N591;
	assign N1066 = N592;
	assign N1148 = ~N592;
	assign N1067 = ~N595;
	assign N1080 = ~N596;
	assign N1092 = ~N597;
	assign N1104 = ~N598;
	assign N2624 = ~( AND3_242_inw1 | N599 );
	assign N7464 = ~( AND3_1945_inw1 | N599 );
	assign N1755 = ~N599;
	assign AND3_1792_inw1 = ~( N6979 & N603 );
	assign AND3_1945_inw1 = ~( N7250 & N603 );
	assign N1758 = ~N603;
	assign N2605 = ~( AND3_223_inw1 | N607 );
	assign N2606 = ~( AND3_224_inw1 | N607 );
	assign N2607 = ~( AND3_225_inw1 | N607 );
	assign N2608 = ~( AND3_226_inw1 | N607 );
	assign N2609 = ~( AND3_227_inw1 | N607 );
	assign N2610 = ~( AND3_228_inw1 | N607 );
	assign N2611 = ~( AND3_229_inw1 | N607 );
	assign N2612 = ~( AND3_230_inw1 | N607 );
	assign N2613 = ~( AND3_231_inw1 | N607 );
	assign N2614 = ~( AND3_232_inw1 | N607 );
	assign N3641 = ~( AND3_600_inw1 | N607 );
	assign N3642 = ~( AND3_601_inw1 | N607 );
	assign N3643 = ~( AND3_602_inw1 | N607 );
	assign N3644 = ~( AND3_603_inw1 | N607 );
	assign N3645 = ~( AND3_604_inw1 | N607 );
	assign N3646 = ~( AND3_605_inw1 | N607 );
	assign N3647 = ~( AND3_606_inw1 | N607 );
	assign N3648 = ~( AND3_607_inw1 | N607 );
	assign N3649 = ~( AND3_608_inw1 | N607 );
	assign N3650 = ~( AND3_609_inw1 | N607 );
	assign N2790 = ~N607;
	assign AND3_1883_inw1 = ~( N7190 & N610 );
	assign AND3_1932_inw1 = ~( N7304 & N610 );
	assign AND3_1934_inw1 = ~( N7282 & N610 );
	assign AND3_1936_inw1 = ~( N7276 & N610 );
	assign AND3_1937_inw1 = ~( N7270 & N610 );
	assign AND3_2052_inw1 = ~( N7549 & N610 );
	assign AND3_2054_inw1 = ~( N7543 & N610 );
	assign AND3_2056_inw1 = ~( N7537 & N610 );
	assign AND3_2058_inw1 = ~( N7531 & N610 );
	assign AND3_2293_inw1 = ~( N8093 & N610 );
	assign N2779 = ~N610;
	assign AND3_1887_inw1 = ~( N7190 & N613 );
	assign AND3_1939_inw1 = ~( N7304 & N613 );
	assign AND3_1941_inw1 = ~( N7282 & N613 );
	assign AND3_1943_inw1 = ~( N7276 & N613 );
	assign AND3_1944_inw1 = ~( N7270 & N613 );
	assign AND3_2050_inw1 = ~( N7549 & N613 );
	assign AND3_2060_inw1 = ~( N7543 & N613 );
	assign AND3_2062_inw1 = ~( N7537 & N613 );
	assign AND3_2064_inw1 = ~( N7531 & N613 );
	assign AND3_2295_inw1 = ~( N8093 & N613 );
	assign N2801 = ~N613;
	assign N2604 = ~( AND3_222_inw1 | N616 );
	assign N2615 = ~( AND3_233_inw1 | N616 );
	assign N2616 = ~( AND3_234_inw1 | N616 );
	assign N2617 = ~( AND3_235_inw1 | N616 );
	assign N2618 = ~( AND3_236_inw1 | N616 );
	assign N2619 = ~( AND3_237_inw1 | N616 );
	assign N2620 = ~( AND3_238_inw1 | N616 );
	assign N2621 = ~( AND3_239_inw1 | N616 );
	assign N2622 = ~( AND3_240_inw1 | N616 );
	assign N2626 = ~( AND3_244_inw1 | N616 );
	assign N3638 = ~( AND3_597_inw1 | N616 );
	assign N3651 = ~( AND3_610_inw1 | N616 );
	assign N3652 = ~( AND3_611_inw1 | N616 );
	assign N3653 = ~( AND3_612_inw1 | N616 );
	assign N3654 = ~( AND3_613_inw1 | N616 );
	assign N3655 = ~( AND3_614_inw1 | N616 );
	assign N3656 = ~( AND3_615_inw1 | N616 );
	assign N3657 = ~( AND3_616_inw1 | N616 );
	assign N3658 = ~( AND3_617_inw1 | N616 );
	assign N3660 = ~( AND3_619_inw1 | N616 );
	assign N2812 = ~N616;
	assign N2625 = ( N619 & N625 );
	assign N8077 = ( N8073 & N619 );
	assign N8078 = ( N8074 & N619 );
	assign AND3_1589_inw1 = ~( N6164 & N619 );
	assign AND3_1803_inw1 = ~( N6932 & N619 );
	assign AND3_1804_inw1 = ~( N6967 & N619 );
	assign AND3_1834_inw1 = ~( N7037 & N619 );
	assign AND3_1835_inw1 = ~( N7034 & N619 );
	assign AND3_1836_inw1 = ~( N7031 & N619 );
	assign AND3_1838_inw1 = ~( N7060 & N619 );
	assign AND3_1839_inw1 = ~( N7057 & N619 );
	assign AND3_1844_inw1 = ~( N7028 & N619 );
	assign AND3_1845_inw1 = ~( N7054 & N619 );
	assign AND3_1958_inw1 = ~( N7245 & N619 );
	assign AND3_1959_inw1 = ~( N7242 & N619 );
	assign AND3_1960_inw1 = ~( N7239 & N619 );
	assign AND3_1961_inw1 = ~( N7236 & N619 );
	assign AND3_1962_inw1 = ~( N7263 & N619 );
	assign AND3_1963_inw1 = ~( N7260 & N619 );
	assign AND3_1964_inw1 = ~( N7257 & N619 );
	assign AND3_1965_inw1 = ~( N7250 & N619 );
	assign AND3_2274_inw1 = ~( N8064 & N619 );
	assign AND3_2275_inw1 = ~( N8061 & N619 );
	assign N3068 = ~N619;
	assign N3659 = ~( AND3_618_inw1 | N625 );
	assign N3661 = ~( AND3_620_inw1 | N625 );
	assign N3781 = ~( AND3_717_inw1 | N625 );
	assign N3782 = ~( AND3_718_inw1 | N625 );
	assign N3783 = ~( AND3_719_inw1 | N625 );
	assign N3784 = ~( AND3_720_inw1 | N625 );
	assign N3785 = ~( AND3_721_inw1 | N625 );
	assign N3786 = ~( AND3_722_inw1 | N625 );
	assign N3787 = ~( AND3_723_inw1 | N625 );
	assign N3788 = ~( AND3_724_inw1 | N625 );
	assign N3800 = ~( AND3_728_inw1 | N625 );
	assign N3801 = ~( AND3_729_inw1 | N625 );
	assign N3802 = ~( AND3_730_inw1 | N625 );
	assign N3803 = ~( AND3_731_inw1 | N625 );
	assign N3804 = ~( AND3_732_inw1 | N625 );
	assign N3805 = ~( AND3_733_inw1 | N625 );
	assign N3806 = ~( AND3_734_inw1 | N625 );
	assign N3807 = ~( AND3_735_inw1 | N625 );
	assign N3808 = ~( AND3_736_inw1 | N625 );
	assign N3809 = ~( AND3_737_inw1 | N625 );
	assign N3063 = ~N625;
	assign N1972 = ~N1146;
	assign N6512 = ( N4310 | N6107 );
	assign g32_inw2 = ~( N5431 & N6107 );
	assign N6817 = ( N6397 | N6664 );
	assign N6106 = ~( AND3_1351_inw1 | N5452 );
	assign N6104 = ~( AND4_1349_inw1 | AND4_1349_inw2 );
	assign N6932 = ~( N6650 & N6806 );
	assign N6650 = ~( N5462 & N2637 );
	assign N4038 = ~( AND3_813_inw1 | N1475 );
	assign N4032 = ~( AND3_807_inw1 | N1475 );
	assign N4033 = ~( AND3_808_inw1 | N1475 );
	assign N4034 = ~( AND3_809_inw1 | N1475 );
	assign N2060 = ~N1150;
	assign N4031 = ( N3828 & N1475 );
	assign N4036 = ( N3829 & N1475 );
	assign N4042 = ( N3831 & N1475 );
	assign N4035 = ~( AND3_810_inw1 | N1475 );
	assign N4037 = ~( AND3_812_inw1 | N1475 );
	assign N4039 = ~( AND3_814_inw1 | N1475 );
	assign N4040 = ~( AND3_815_inw1 | N1475 );
	assign N2623 = ~N1475;
	assign N3829 = ( N3740 | N2971 );
	assign N5346 = ( N3921 | N5119 );
	assign g28_inw2 = ~( N5264 & N5119 );
	assign N6844 = ( N6427 | N6693 );
	assign N6163 = ~( AND3_1400_inw1 | N5606 );
	assign N6161 = ~( AND4_1398_inw1 | AND4_1398_inw2 );
	assign N6164 = ~( N5616 & N5955 );
	assign N5616 = ~( N4405 & N2715 );
	assign N3831 = ( N3738 | N2969 );
	assign N3828 = ( N3739 | N2970 );
	assign N8096 = ( N8090 | N3072 );
	assign N8093 = ( N8089 | N3071 );
	assign N6979 = ( N6879 | N6880 );
	assign N6879 = ( N4357 & N6478 );
	assign N1149 = ~N1042;
	assign N8127 = ~N8125;
	assign N8128 = ~N8126;
	assign N3893 = ( N3689 | N2876 );
	assign OR3_836_inw1 = ~( N3761 | N3982 );
	assign N4183 = ( N3758 | N3980 );
	assign N4264 = ~( N4024 & N3823 );
	assign N3980 = ~( AND3_790_inw1 | N3753 );
	assign OR3_627_inw1 = ~( N2835 | N3405 );
	assign OR3_709_inw1 = ~( N3027_key | N3508_key );
	assign N3887 = ( N3688 | N2875 );
	assign N3664 = ( N2831 | N3401 );
	assign N3763 = ( N3023_key | N3504 );
	assign N3405 = ( N1080 & N2823 );
	assign N3401 = ~( AND3_495_inw1 | N2823 );
	assign N3504 = ~( AND3_547_inw1_key | N2823 );
	assign OR3_628_inw1 = ~( N2836 | N3406 );
	assign OR3_710_inw1 = ~( N3028_key | N3509_key );
	assign N3881 = ( N3687 | N2874 );
	assign N3665 = ( N2832 | N3402 );
	assign N3764 = ( N3024_key | N3505 );
	assign N3824 = ~( N3609 & N3610 );
	assign N3406 = ( N1080 & N2825 );
	assign N3402 = ~( AND3_496_inw1 | N2825 );
	assign N3505 = ~( AND3_548_inw1_key | N2825 );
	assign OR3_629_inw1 = ~( N2837 | N3407 );
	assign OR3_711_inw1 = ~( N3029_key | N3510_key );
	assign N3873 = ( N3686 | N2873 );
	assign N3666 = ( N2833 | N3403 );
	assign N3765 = ( N3025_key | N3506 );
	assign N3407 = ( N1080 & N2827 );
	assign N3403 = ~( AND3_497_inw1 | N2827 );
	assign N3506 = ~( AND3_549_inw1_key | N2827 );
	assign OR3_630_inw1 = ~( N2838 | N3408 );
	assign OR3_712_inw1 = ~( N3030_key | N3511_key );
	assign N3867 = ( N3685 | N2872 );
	assign N3667 = ( N2834 | N3404 );
	assign N3766 = ( N3026_key | N3507 );
	assign N3797 = ~( N3562 & N3563 );
	assign N3408 = ( N1080 & N2829 );
	assign N3404 = ~( AND3_498_inw1 | N2829 );
	assign N3507 = ~( AND3_550_inw1_key | N2829 );
	assign N3705 = ( N2910 | N3447 );
	assign OR3_653_inw1 = ~( N2911 | N3448 );
	assign OR3_654_inw1 = ~( N2912 | N3449 );
	assign OR3_666_inw1 = ~( N2938_key | N3463_key );
	assign OR3_667_inw1 = ~( N2939_key | N3464_key );
	assign OR3_668_inw1 = ~( N2940_key | N3465_key );
	assign OR3_669_inw1 = ~( N2941_key | N3466_key );
	assign OR3_687_inw1 = ~( N2983 | N3485 );
	assign OR3_688_inw1 = ~( N2985 | N3486 );
	assign OR3_689_inw1 = ~( N2986 | N3487 );
	assign N3816 = ( N3482 & N2984 );
	assign g49_inw2 = ~( n_330 & n_331 );
	assign N3700 = ( N2907 | N3444 );
	assign N3482 = ~N2980;
	assign N3757 = ( N3013 | N3502 );
	assign N3445 = ~( AND3_512_inw1 | N2903 );
	assign N3446 = ~( AND3_513_inw1 | N2905 );
	assign N3459 = ~( AND3_524_inw1_key | N2839 );
	assign N3460 = ~( AND3_525_inw1_key | N2841 );
	assign N3461 = ~( AND3_526_inw1_key | N2843 );
	assign N3462 = ~( AND3_527_inw1_key | N2845 );
	assign N3481 = ~( AND3_532_inw1 | N1660 );
	assign N3483 = ~( AND3_534_inw1 | N2915 );
	assign N3484 = ~( AND3_535_inw1 | N2917 );
	assign OR3_635_inw1 = ~( N2851 | N3413 );
	assign N3861 = ( N3684 | N2871 );
	assign N3672 = ( N2847 | N3409 );
	assign N3715 = ( N2934_key | N3459 );
	assign N3413 = ( N1080 & N2839 );
	assign N3409 = ~( AND3_503_inw1 | N2839 );
	assign OR3_636_inw1 = ~( N2852 | N3414 );
	assign N3855 = ( N3683 | N2870 );
	assign N3673 = ( N2848 | N3410 );
	assign N3716 = ( N2935_key | N3460 );
	assign N3793 = ~( N3560 & N3561 );
	assign N3414 = ( N1080 & N2841 );
	assign N3410 = ~( AND3_504_inw1 | N2841 );
	assign OR3_637_inw1 = ~( N2853 | N3415 );
	assign N3849 = ( N3682 | N2869 );
	assign N3674 = ( N2849 | N3411 );
	assign N3717 = ( N2936_key | N3461 );
	assign N3415 = ( N1080 & N2843 );
	assign N3411 = ~( AND3_505_inw1 | N2843 );
	assign OR3_638_inw1 = ~( N2854 | N3416 );
	assign N3842 = ( N3681 | N2868 );
	assign N3675 = ( N2850 | N3412 );
	assign N3718 = ( N2937_key | N3462 );
	assign N3789 = ~( N3558 & N3559 );
	assign N3416 = ( N1080 & N2845 );
	assign N3412 = ~( AND3_506_inw1 | N2845 );
	assign N4011 = ( N3680_key | N2867_key );
	assign N3968 = ( N3731 | N2963 );
	assign N3810 = ~( N3607 & N3608 );
	assign N3962 = ( N3730 | N2962 );
	assign N3956 = ( N3729 | N2961 );
	assign N3701 = ( N2908 | N3445 );
	assign N3813 = ~( N3605 & N3606 );
	assign N3948 = ( N3728 | N2960 );
	assign N3702 = ( N2909 | N3446 );
	assign OR3_659_inw1 = ~( N2923 | N3453 );
	assign N3942 = ( N3727 | N2959 );
	assign N3708 = ( N2919 | N3450 );
	assign N3742 = ( N2979 | N3481 );
	assign N5147 = ~( N4953 | N4196 );
	assign N5148 = ~( N4954 | N4955 );
	assign N3453 = ( N1080 & N1660 );
	assign N3450 = ~( AND3_517_inw1 | N1660 );
	assign N4196 = ~( AND3_840_inw1 | N1660 );
	assign N4955 = ~( AND3_1005_inw1 | N1660 );
	assign N4008 = ( N3723_key | N2954_key );
	assign N3921 = ( N3724 | N2955 );
	assign N3927 = ( N3725 | N2956 );
	assign N3933 = ( N3726 | N2957 );
	assign N3732 = ( N2942 | N2958 );
	assign OR3_660_inw1 = ~( N2924 | N3454 );
	assign N3709 = ( N2921 | N3451 );
	assign N3743 = ( N2981 | N3483 );
	assign N3775 = ~( N3514 & N3515 );
	assign N3454 = ( N1080 & N2915 );
	assign N3451 = ~( AND3_518_inw1 | N2915 );
	assign OR3_661_inw1 = ~( N2925 | N3455 );
	assign N3710 = ( N2922 | N3452 );
	assign N3744 = ( N2982 | N3484 );
	assign N3455 = ( N1080 & N2917 );
	assign N3452 = ~( AND3_519_inw1 | N2917 );
	assign N3771 = ~( N3512 & N3513 );
	assign N6105 = ( N5452 & N4310 );
	assign N6103 = ~( AND3_1348_inw1 | N4310 );
	assign AND4_1345_inw2 = ~( N4310 & N5431 );
	assign N6990 = ~( N4310 & N6895 );
	assign N5728 = ~N4310;
	assign g12_inw1 = ~( N5424 & N4310 );
	assign N5462 = ~( N5250 & N5086 );
	assign N6987 = ~( N4608_key & N6889 );
	assign N5176 = ~N4608_key;
	assign N5086 = ~( N3842 & N2636 );
	assign N4109 = ( N3841 & N3679 );
	assign N4198 = ( N3920 & N3722_key );
	assign N2061 = ~N1151;
	assign N6094 = ( N5424 & N4298 );
	assign NOR4_1525_inw1 = ~( N4298 | N6098 );
	assign n_316 = ( N4298 | N6098 );
	assign N5431 = ~( N5247 & N5080 );
	assign N5080 = ~( N3861 & N2633 );
	assign N4100 = ( N3838 & N3676 );
	assign N4234 = ( N3917 & N3719_key );
	assign N6098 = ( N5431 & N4301 );
	assign N6095 = ~( AND3_1340_inw1 | N4301 );
	assign NOR3_1524_inw1 = ~( N4301 | N6102 );
	assign OR4_1517_inw1 = ~( N4301 | N6102 );
	assign OR4_1522_inw1 = ~( N4301 | N6102 );
	assign N5441 = ~( N5248 & N5082 );
	assign N5082 = ~( N3855 & N2634 );
	assign N4103 = ( N3839 & N3677 );
	assign N4225 = ( N3918 & N3720_key );
	assign N6102 = ( N4305 & N5441 );
	assign AND3_1344_inw1 = ~( N5441 & N4305 );
	assign AND4_1341_inw2 = ~( N4305 & N5431 );
	assign N6419 = ( N4305 | N6105 );
	assign OR3_1518_inw1 = ~( N4305 | N6105 );
	assign N5452 = ~( N5249 & N5084 );
	assign N5084 = ~( N3849 & N2635 );
	assign N4106 = ( N3840 & N3678 );
	assign N4228 = ( N3919 & N3721_key );
	assign N6088 = ( N5407 & N4290 );
	assign AND3_1331_inw1 = ~( N5407 & N4290 );
	assign AND4_1322_inw2 = ~( N4290 & N5396 );
	assign N6816 = ~( N4290 & N6661 );
	assign N7153 = ~( N4290 & N6411 );
	assign N5469 = ~N4290;
	assign N5418 = ~( N5245 & N5076 );
	assign N6815 = ~( N4575 & N6661 );
	assign N7152 = ~( N4575 & N7072 );
	assign N5087 = ~N4575;
	assign N5076 = ~( N3873 & N2631 );
	assign N4094 = ( N3836 & N3670 );
	assign N4240 = ( N3990 & N3769_key );
	assign n_306 = ( N4297 | N6094 );
	assign N5424 = ~( N5246 & N5078 );
	assign N5078 = ~( N3867 & N2632 );
	assign N4097 = ( N3837 & N3671 );
	assign N4231 = ( N3991 & N3770_key );
	assign OR4_1486_inw1 = ~( N4268 | N6071 );
	assign N5389 = ~( N5242 & N5070 );
	assign N5070 = ~( N3893 & N2628 );
	assign N4939 = ( N4515 & N4185 );
	assign N6071 = ( N5389 & N4280 );
	assign NOR3_1513_inw1 = ~( N4280 | N6083 );
	assign OR4_1512_inw1 = ~( N4280 | N6083 );
	assign N5396 = ~( N5243 & N5072 );
	assign N5072 = ~( N3887 & N2629 );
	assign N4088 = ( N3834 & N3668 );
	assign N4243 = ( N3988 & N3767 );
	assign N6083 = ( N5396 & N4284 );
	assign N6072 = ~( AND3_1321_inw1 | N4284 );
	assign N6494 = ~( N4284 | N6088 );
	assign OR3_1514_inw1 = ~( N4284 | N6088 );
	assign N5407 = ~( N5244 & N5074 );
	assign N5074 = ~( N3881 & N2630 );
	assign N4091 = ( N3835 & N3669 );
	assign N4237 = ( N3989 & N3768 );
	assign N5117 = ( N4364 & N4379 );
	assign N5066 = ~( AND3_1046_inw1 | N4379 );
	assign N6575 = ~( N4379 | N6146 );
	assign OR3_1528_inw1 = ~( N4379 | N6146 );
	assign N5562 = ~( N5261 & N5107 );
	assign N5107 = ~( N3956 & N2709 );
	assign N4144 = ( N3908 & N3703 );
	assign N6146 = ( N5562 & N4385 );
	assign AND3_1382_inw1 = ~( N5562 & N4385 );
	assign AND4_1323_inw2 = ~( N4385 & N4364 );
	assign N6843 = ~( N4385 & N6690 );
	assign N7159 = ~( N4385 & N6437 );
	assign N5622 = ~N4385;
	assign N5573 = ~( N5262 & N5109 );
	assign N6842 = ~( N4627 & N6690 );
	assign N7158 = ~( N4627 & N7084 );
	assign N5120 = ~N4627;
	assign N5109 = ~( N3948 & N2710 );
	assign N4147 = ( N3909 & N3704 );
	assign n_308 = ( N4392 | N6152 );
	assign N5579 = ~( N5263 & N5111 );
	assign N5111 = ~( N3942 & N2711 );
	assign N4153 = ( N3914 & N3711 );
	assign N4252 = ( N3975 & N3745 );
	assign N2920 = ~N2349;
	assign N6152 = ( N5579 & N4067 );
	assign NOR4_1538_inw1 = ~( N4067 | N5954 );
	assign n_314 = ( N4067 | N5954 );
	assign N5264 = ~( N5112 & N4856 );
	assign N4856 = ~( N3732 & N2712 );
	assign N3456 = ( N2920 & N2350 );
	assign N5954 = ( N5264 & N4396 );
	assign N6153 = ~( AND3_1390_inw1 | N4396 );
	assign NOR3_1537_inw1 = ~( N4396 | N6159 );
	assign OR4_1531_inw1 = ~( N4396 | N6159 );
	assign OR4_1535_inw1 = ~( N4396 | N6159 );
	assign N5595 = ~( N5274 & N5114 );
	assign N5114 = ~( N3933 & N2713 );
	assign N4156 = ( N3915 & N3712 );
	assign N4246 = ( N3976 & N3746 );
	assign N6159 = ( N4400 & N5595 );
	assign AND3_1393_inw1 = ~( N5595 & N4400 );
	assign AND4_1391_inw2 = ~( N4400 & N5264 );
	assign N6445 = ( N4400 | N6162 );
	assign OR3_1532_inw1 = ~( N4400 | N6162 );
	assign N5606 = ~( N5275 & N5116 );
	assign N5116 = ~( N3927 & N2714 );
	assign N4159 = ( N3916 & N3713 );
	assign N4249 = ( N3977 & N3747 );
	assign N1143 = N1137;
	assign N1142 = N1137;
	assign N2584 = N1141;
	assign g49_inw1 = ~( n_328 & n_329 );
	assign N8045 = ( N8043 | N8041 );
	assign OR4_2241_inw2 = ~( N7990 | N7991 );
	assign N8043 = ( N8040 & N1157 );
	assign N7988 = ~( AND3_2227_inw1 | N1157 );
	assign N7989 = ~( AND3_2228_inw1 | N1157 );
	assign N7338 = ~( AND3_1879_inw1 | N2664 );
	assign N7434 = ~( AND3_1915_inw1 | N2664 );
	assign N7436 = ~( AND3_1917_inw1 | N2664 );
	assign N7438 = ~( AND3_1919_inw1 | N2664 );
	assign N7440 = ~( AND3_1921_inw1 | N2664 );
	assign N7667 = ~( AND3_2034_inw1 | N2664 );
	assign N7669 = ~( AND3_2036_inw1 | N2664 );
	assign N7671 = ~( AND3_2038_inw1 | N2664 );
	assign N7673 = ~( AND3_2040_inw1 | N2664 );
	assign N8118 = ~( AND3_2297_inw1 | N2664 );
	assign AND3_1743_inw1 = ~( N6866 & N2653 );
	assign AND3_1880_inw1 = ~( N7198 & N2653 );
	assign AND3_1914_inw1 = ~( N7310 & N2653 );
	assign AND3_1918_inw1 = ~( N7288 & N2653 );
	assign AND3_1920_inw1 = ~( N7294 & N2653 );
	assign AND3_2033_inw1 = ~( N7555 & N2653 );
	assign AND3_2035_inw1 = ~( N7561 & N2653 );
	assign AND3_2037_inw1 = ~( N7567 & N2653 );
	assign AND3_2039_inw1 = ~( N7573 & N2653 );
	assign AND3_2296_inw1 = ~( N8096 & N2653 );
	assign OR4_1974_inw2 = ~( N3616 | N2585 );
	assign OR4_2088_inw2 = ~( N3617 | N2586 );
	assign OR4_2089_inw2 = ~( N3618 | N2587 );
	assign OR4_2090_inw2 = ~( N3619 | N2588 );
	assign OR4_2091_inw2 = ~( N3620 | N2589 );
	assign OR4_1916_inw2 = ~( N3621 | N2591 );
	assign OR4_1976_inw2 = ~( N3622 | N2592 );
	assign OR4_1977_inw2 = ~( N3623 | N2593 );
	assign OR4_1978_inw2 = ~( N3624 | N2594 );
	assign OR4_2300_inw2 = ~( N3662 | N2703 );
	assign N7011 = ~( AND3_1743_inw1 | N2664 );
	assign N7339 = ~( AND3_1880_inw1 | N2664 );
	assign N7433 = ~( AND3_1914_inw1 | N2664 );
	assign N7437 = ~( AND3_1918_inw1 | N2664 );
	assign N7439 = ~( AND3_1920_inw1 | N2664 );
	assign N7666 = ~( AND3_2033_inw1 | N2664 );
	assign N7668 = ~( AND3_2035_inw1 | N2664 );
	assign N7670 = ~( AND3_2037_inw1 | N2664 );
	assign N7672 = ~( AND3_2039_inw1 | N2664 );
	assign N8117 = ~( AND3_2296_inw1 | N2664 );
	assign N7340 = ~( AND3_1881_inw1 | N2739 );
	assign N7442 = ~( AND3_1923_inw1 | N2739 );
	assign N7444 = ~( AND3_1925_inw1 | N2739 );
	assign N7446 = ~( AND3_1927_inw1 | N2739 );
	assign N7448 = ~( AND3_1929_inw1 | N2739 );
	assign N7675 = ~( AND3_2042_inw1 | N2739 );
	assign N7677 = ~( AND3_2044_inw1 | N2739 );
	assign N7679 = ~( AND3_2046_inw1 | N2739 );
	assign N7681 = ~( AND3_2048_inw1 | N2739 );
	assign N8120 = ~( AND3_2299_inw1 | N2739 );
	assign AND3_1744_inw1 = ~( N6866 & N2728 );
	assign AND3_1882_inw1 = ~( N7198 & N2728 );
	assign AND3_1922_inw1 = ~( N7310 & N2728 );
	assign AND3_1926_inw1 = ~( N7288 & N2728 );
	assign AND3_1928_inw1 = ~( N7294 & N2728 );
	assign AND3_2041_inw1 = ~( N7555 & N2728 );
	assign AND3_2043_inw1 = ~( N7561 & N2728 );
	assign AND3_2045_inw1 = ~( N7567 & N2728 );
	assign AND3_2047_inw1 = ~( N7573 & N2728 );
	assign AND3_2298_inw1 = ~( N8096 & N2728 );
	assign OR4_1979_inw2 = ~( N3627 | N2595 );
	assign OR4_2092_inw2 = ~( N3628 | N2596 );
	assign OR4_2093_inw2 = ~( N3629 | N2597 );
	assign OR4_2094_inw2 = ~( N3630 | N2598 );
	assign OR4_2095_inw2 = ~( N3631 | N2599 );
	assign OR4_1924_inw2 = ~( N3632 | N2600 );
	assign OR4_1981_inw2 = ~( N3633 | N2601 );
	assign OR4_1982_inw2 = ~( N3634 | N2602 );
	assign OR4_1983_inw2 = ~( N3635 | N2603 );
	assign OR4_2301_inw2 = ~( N3663 | N2778 );
	assign N7012 = ~( AND3_1744_inw1 | N2739 );
	assign N7341 = ~( AND3_1882_inw1 | N2739 );
	assign N7441 = ~( AND3_1922_inw1 | N2739 );
	assign N7445 = ~( AND3_1926_inw1 | N2739 );
	assign N7447 = ~( AND3_1928_inw1 | N2739 );
	assign N7674 = ~( AND3_2041_inw1 | N2739 );
	assign N7676 = ~( AND3_2043_inw1 | N2739 );
	assign N7678 = ~( AND3_2045_inw1 | N2739 );
	assign N7680 = ~( AND3_2047_inw1 | N2739 );
	assign N8119 = ~( AND3_2298_inw1 | N2739 );
	assign N8048 = ( N8044 | N8035 );
	assign OR4_2242_inw2 = ~( N7996 | N7997 );
	assign N8044 = ( N8042 & N1219 );
	assign N7994 = ~( AND3_2233_inw1 | N1219 );
	assign N7995 = ~( AND3_2234_inw1 | N1219 );
	assign OR4_873_inw2 = ~( N3614 | N3615 );
	assign OR4_874_inw2 = ~( N3614 | N3615 );
	assign OR4_876_inw2 = ~( N3614 | N3615 );
	assign OR4_877_inw2 = ~( N3614 | N3615 );
	assign N3614 = ( N1588 & N2623 );
	assign OR4_1992_inw2 = ~( N2624 | N7464 );
	assign N4741 = ~( AND3_995_inw1 | N1755 );
	assign N7114 = ~( AND3_1792_inw1 | N1755 );
	assign AND3_995_inw1 = ~( N3705 & N1758 );
	assign OR4_1930_inw2 = ~( N3641 | N2605 );
	assign OR4_2097_inw2 = ~( N3642 | N2606 );
	assign OR4_2098_inw2 = ~( N3643 | N2607 );
	assign OR4_2099_inw2 = ~( N3644 | N2608 );
	assign OR4_2100_inw2 = ~( N3645 | N2609 );
	assign OR4_1984_inw2 = ~( N3646 | N2610 );
	assign OR4_1985_inw2 = ~( N3647 | N2611 );
	assign OR4_1986_inw2 = ~( N3648 | N2612 );
	assign OR4_1987_inw2 = ~( N3649 | N2613 );
	assign OR4_2302_inw2 = ~( N3650 | N2614 );
	assign N7013 = ~( AND3_1745_inw1 | N2790 );
	assign N7342 = ~( AND3_1883_inw1 | N2790 );
	assign N7349 = ~( AND3_1884_inw1 | N2790 );
	assign N7450 = ~( AND3_1931_inw1 | N2790 );
	assign N7451 = ~( AND3_1932_inw1 | N2790 );
	assign N7452 = ~( AND3_1933_inw1 | N2790 );
	assign N7453 = ~( AND3_1934_inw1 | N2790 );
	assign N7454 = ~( AND3_1935_inw1 | N2790 );
	assign N7455 = ~( AND3_1936_inw1 | N2790 );
	assign N7456 = ~( AND3_1937_inw1 | N2790 );
	assign N7684 = ~( AND3_2051_inw1 | N2790 );
	assign N7685 = ~( AND3_2052_inw1 | N2790 );
	assign N7686 = ~( AND3_2053_inw1 | N2790 );
	assign N7687 = ~( AND3_2054_inw1 | N2790 );
	assign N7688 = ~( AND3_2055_inw1 | N2790 );
	assign N7689 = ~( AND3_2056_inw1 | N2790 );
	assign N7690 = ~( AND3_2057_inw1 | N2790 );
	assign N7691 = ~( AND3_2058_inw1 | N2790 );
	assign N8113 = ~( AND3_2292_inw1 | N2790 );
	assign N8114 = ~( AND3_2293_inw1 | N2790 );
	assign AND3_1745_inw1 = ~( N6866 & N2779 );
	assign AND3_1884_inw1 = ~( N7198 & N2779 );
	assign AND3_1931_inw1 = ~( N7310 & N2779 );
	assign AND3_1933_inw1 = ~( N7294 & N2779 );
	assign AND3_1935_inw1 = ~( N7288 & N2779 );
	assign AND3_2051_inw1 = ~( N7573 & N2779 );
	assign AND3_2053_inw1 = ~( N7567 & N2779 );
	assign AND3_2055_inw1 = ~( N7561 & N2779 );
	assign AND3_2057_inw1 = ~( N7555 & N2779 );
	assign AND3_2292_inw1 = ~( N8096 & N2779 );
	assign N7364 = ~( AND3_1887_inw1 | N2812 );
	assign N7458 = ~( AND3_1939_inw1 | N2812 );
	assign N7460 = ~( AND3_1941_inw1 | N2812 );
	assign N7462 = ~( AND3_1943_inw1 | N2812 );
	assign N7463 = ~( AND3_1944_inw1 | N2812 );
	assign N7683 = ~( AND3_2050_inw1 | N2812 );
	assign N7693 = ~( AND3_2060_inw1 | N2812 );
	assign N7695 = ~( AND3_2062_inw1 | N2812 );
	assign N7697 = ~( AND3_2064_inw1 | N2812 );
	assign N8116 = ~( AND3_2295_inw1 | N2812 );
	assign AND3_1747_inw1 = ~( N6866 & N2801 );
	assign AND3_1885_inw1 = ~( N7198 & N2801 );
	assign AND3_1938_inw1 = ~( N7310 & N2801 );
	assign AND3_1940_inw1 = ~( N7294 & N2801 );
	assign AND3_1942_inw1 = ~( N7288 & N2801 );
	assign AND3_2049_inw1 = ~( N7573 & N2801 );
	assign AND3_2059_inw1 = ~( N7567 & N2801 );
	assign AND3_2061_inw1 = ~( N7561 & N2801 );
	assign AND3_2063_inw1 = ~( N7555 & N2801 );
	assign AND3_2294_inw1 = ~( N8096 & N2801 );
	assign OR4_2096_inw2 = ~( N3638 | N2604 );
	assign OR4_2101_inw2 = ~( N3651 | N2615 );
	assign OR4_2102_inw2 = ~( N3652 | N2616 );
	assign OR4_2103_inw2 = ~( N3653 | N2617 );
	assign OR4_1988_inw2 = ~( N3654 | N2618 );
	assign OR4_1989_inw2 = ~( N3655 | N2619 );
	assign OR4_1990_inw2 = ~( N3656 | N2620 );
	assign OR4_1991_inw2 = ~( N3657 | N2621 );
	assign OR4_2303_inw2 = ~( N3658 | N2622 );
	assign OR4_1950_inw2 = ~( N3660 | N2626 );
	assign N7016 = ~( AND3_1747_inw1 | N2812 );
	assign N7357 = ~( AND3_1885_inw1 | N2812 );
	assign N7457 = ~( AND3_1938_inw1 | N2812 );
	assign N7459 = ~( AND3_1940_inw1 | N2812 );
	assign N7461 = ~( AND3_1942_inw1 | N2812 );
	assign N7682 = ~( AND3_2049_inw1 | N2812 );
	assign N7692 = ~( AND3_2059_inw1 | N2812 );
	assign N7694 = ~( AND3_2061_inw1 | N2812 );
	assign N7696 = ~( AND3_2063_inw1 | N2812 );
	assign N8115 = ~( AND3_2294_inw1 | N2812 );
	assign OR4_2278_inw2 = ~( N3659 | N2625 );
	assign OR4_2279_inw2 = ~( N3661 | N2625 );
	assign N8079 = ( N7530 | N8077 );
	assign N8082 = ( N7479 | N8078 );
	assign N6718 = ~( AND3_1589_inw1 | N3063 );
	assign N7146 = ~( AND3_1803_inw1 | N3063 );
	assign N7147 = ~( AND3_1804_inw1 | N3063 );
	assign N7187 = ~( AND3_1834_inw1 | N3063 );
	assign N7188 = ~( AND3_1835_inw1 | N3063 );
	assign N7189 = ~( AND3_1836_inw1 | N3063 );
	assign N7196 = ~( AND3_1838_inw1 | N3063 );
	assign N7197 = ~( AND3_1839_inw1 | N3063 );
	assign N7207 = ~( AND3_1844_inw1 | N3063 );
	assign N7208 = ~( AND3_1845_inw1 | N3063 );
	assign N7481 = ~( AND3_1958_inw1 | N3063 );
	assign N7482 = ~( AND3_1959_inw1 | N3063 );
	assign N7483 = ~( AND3_1960_inw1 | N3063 );
	assign N7484 = ~( AND3_1961_inw1 | N3063 );
	assign N7485 = ~( AND3_1962_inw1 | N3063 );
	assign N7486 = ~( AND3_1963_inw1 | N3063 );
	assign N7487 = ~( AND3_1964_inw1 | N3063 );
	assign N7488 = ~( AND3_1965_inw1 | N3063 );
	assign N8071 = ~( AND3_2274_inw1 | N3063 );
	assign N8072 = ~( AND3_2275_inw1 | N3063 );
	assign N7479 = ( N7301_key & N3068 );
	assign N7530 = ( N7402_key & N3068 );
	assign AND3_800_inw1 = ~( N3456 & N3068 );
	assign AND3_841_inw1 = ~( N3987 & N3068 );
	assign AND3_923_inw1 = ~( N3911 & N3068 );
	assign AND3_1006_inw1 = ~( N4109 & N3068 );
	assign AND3_1007_inw1 = ~( N4106 & N3068 );
	assign AND3_1008_inw1 = ~( N4103 & N3068 );
	assign AND3_1009_inw1 = ~( N4100 & N3068 );
	assign AND3_1010_inw1 = ~( N4159 & N3068 );
	assign AND3_1011_inw1 = ~( N4156 & N3068 );
	assign AND3_1024_inw1 = ~( N4097 & N3068 );
	assign AND3_1025_inw1 = ~( N4094 & N3068 );
	assign AND3_1026_inw1 = ~( N4091 & N3068 );
	assign AND3_1027_inw1 = ~( N4088 & N3068 );
	assign AND3_1028_inw1 = ~( N4153 & N3068 );
	assign AND3_1029_inw1 = ~( N4147 & N3068 );
	assign AND3_1030_inw1 = ~( N4144 & N3068 );
	assign AND3_1031_inw1 = ~( N3705 & N3068 );
	assign AND3_1139_inw1 = ~( N4939 & N3068 );
	assign AND3_1993_inw1 = ~( N7468 & N3068 );
	assign AND3_2029_inw1 = ~( N7529 & N3068 );
	assign N7190 = ~( OR3_1837_inw1 & N3781 );
	assign N7270 = ~( OR3_1867_inw1 & N3782 );
	assign N7276 = ~( OR3_1868_inw1 & N3783 );
	assign N7282 = ~( OR3_1869_inw1 & N3784 );
	assign N6866 = ~( OR3_1670_inw1 & N3785 );
	assign N7198 = ~( OR3_1840_inw1 & N3786 );
	assign N7288 = ~( OR3_1870_inw1 & N3787 );
	assign N7294 = ~( OR3_1871_inw1 & N3788 );
	assign N7304 = ~( OR3_1874_inw1 & N3800 );
	assign N7531 = ~( OR3_1998_inw1 & N3801 );
	assign N7537 = ~( OR3_1999_inw1 & N3802 );
	assign N7543 = ~( OR3_2000_inw1 & N3803 );
	assign N7549 = ~( OR3_2001_inw1 & N3804 );
	assign N7310 = ~( OR3_1875_inw1 & N3805 );
	assign N7555 = ~( OR3_2002_inw1 & N3806 );
	assign N7561 = ~( OR3_2003_inw1 & N3807 );
	assign N7567 = ~( OR3_2004_inw1 & N3808 );
	assign N7573 = ~( OR3_2005_inw1 & N3809 );
	assign N8089 = ( N8079 & N3063 );
	assign N8090 = ( N8082 & N3063 );
	assign N3998 = ~( AND3_800_inw1 | N3063 );
	assign N4197 = ~( AND3_841_inw1 | N3063 );
	assign N4547 = ~( AND3_923_inw1 | N3063 );
	assign N4956 = ~( AND3_1006_inw1 | N3063 );
	assign N4957 = ~( AND3_1007_inw1 | N3063 );
	assign N4958 = ~( AND3_1008_inw1 | N3063 );
	assign N4959 = ~( AND3_1009_inw1 | N3063 );
	assign N4960 = ~( AND3_1010_inw1 | N3063 );
	assign N4961 = ~( AND3_1011_inw1 | N3063 );
	assign N4980 = ~( AND3_1024_inw1 | N3063 );
	assign N4981 = ~( AND3_1025_inw1 | N3063 );
	assign N4982 = ~( AND3_1026_inw1 | N3063 );
	assign N4983 = ~( AND3_1027_inw1 | N3063 );
	assign N4984 = ~( AND3_1028_inw1 | N3063 );
	assign N4985 = ~( AND3_1029_inw1 | N3063 );
	assign N4986 = ~( AND3_1030_inw1 | N3063 );
	assign N4987 = ~( AND3_1031_inw1 | N3063 );
	assign N5165 = ~( AND3_1139_inw1 | N3063 );
	assign N7526 = ~( AND3_1993_inw1 | N3063 );
	assign N7636 = ~( AND3_2029_inw1 | N3063 );
	assign N6830 = ~( N6512 & N6672 );
	assign N6829 = ~N6512;
	assign N6101 = ~( g32_inw1 | g32_inw2 );
	assign N7040 = ( N6817 & N6079 );
	assign N7125 = ( N6817 & N7018 );
	assign N7126 = ( N6817 & N7020 );
	assign N7127 = ( N6817 & N7022 );
	assign N7023 = ~N6817;
	assign N6508 = ~( OR3_1518_inw1 & N6106 );
	assign OR4_1517_inw2 = ~( N6103 | N6104 );
	assign g33_inw1 = ~( N6932 | N7037 );
	assign OR4_876_inw1 = ~( N4037 | N4038 );
	assign OR4_873_inw1 = ~( N4032 | N4033 );
	assign OR4_874_inw1 = ~( N4034 | N4035 );
	assign N4272 = ~N4031;
	assign N4275 = ~N4036;
	assign N4279 = ~N4042;
	assign OR4_877_inw1 = ~( N4039 | N4040 );
	assign N6856 = ~( N5346 & N6700 );
	assign N5956 = ~N5346;
	assign N6158 = ~( g28_inw1 | g28_inw2 );
	assign N7064 = ( N6844 & N6139 );
	assign N7139 = ( N6844 & N7044 );
	assign N7140 = ( N6844 & N7046 );
	assign N7141 = ( N6844 & N7048 );
	assign N7049 = ~N6844;
	assign N6587 = ~( OR3_1532_inw1 & N6163 );
	assign OR4_1531_inw2 = ~( N6160 | N6161 );
	assign g38_inw1 = ~( N6164 | N6967 );
	assign N7624 = ( N6979 & N7489 );
	assign N7489 = ~( N6979 & N7250 );
	assign N7626 = ( N1149 & N7525 );
	assign N5145 = ~( N3893 & N4523 );
	assign N5069 = ~N3893;
	assign N4515 = ~N4183;
	assign N5059 = ~( N4264 & N4267 );
	assign N5058 = ~N4264;
	assign N5310 = ~( N3887 & N5073 );
	assign N5071 = ~N3887;
	assign N3834 = ~N3664;
	assign N3988 = ~N3763;
	assign N5309 = ~( N3881 & N5071 );
	assign N5073 = ~N3881;
	assign N3835 = ~N3665;
	assign N3989 = ~N3764;
	assign N5239 = ~( N3824 & N5058 );
	assign N4267 = ~N3824;
	assign N5308 = ~( N3873 & N5077 );
	assign N5075 = ~N3873;
	assign N3836 = ~N3666;
	assign N3990 = ~N3765;
	assign N5307 = ~( N3867 & N5075 );
	assign N5077 = ~N3867;
	assign N3837 = ~N3667;
	assign N3991 = ~N3766;
	assign N4978 = ~( AND3_1022_inw1 | N3797 );
	assign N4979 = ~( AND3_1023_inw1 | N3797 );
	assign N4976 = ~N3797;
	assign N5057 = ~( N3705 & N3700 );
	assign N4027 = ~N3705;
	assign N5162 = ~( N3816 & N4974 );
	assign N4199 = ~N3816;
	assign N7703 = ~( g49_inw1 | g49_inw2 );
	assign AND4_1041_inw2 = ~( N3700 & N4027 );
	assign N3911 = ~N3700;
	assign N5240 = ~( AND3_1175_inw1 | N3757 );
	assign AND3_1508_inw1 = ~( N5324 & N3757 );
	assign AND3_1593_inw1 = ~( N3757 & N6028 );
	assign N3987 = ~N3757;
	assign N5370 = ~( N3861 & N5081 );
	assign N5079 = ~N3861;
	assign N3838 = ~N3672;
	assign N3917 = ~N3715;
	assign N5369 = ~( N3855 & N5079 );
	assign N5081 = ~N3855;
	assign N3839 = ~N3673;
	assign N3918 = ~N3716;
	assign AND3_1022_inw1 = ~( N3793 & N3789 );
	assign AND3_1137_inw1 = ~( N4200 & N3793 );
	assign N4203 = ~N3793;
	assign N5368 = ~( N3849 & N5085 );
	assign N5083 = ~N3849;
	assign N3840 = ~N3674;
	assign N3919 = ~N3717;
	assign N5367 = ~( N3842 & N5083 );
	assign N5085 = ~N3842;
	assign N3841 = ~N3675;
	assign N3920 = ~N3718;
	assign AND3_1138_inw1 = ~( N3789 & N4203 );
	assign N4200 = ~N3789;
	assign N5311 = ~( N4011_key & N5069 );
	assign N4523 = ~N4011_key;
	assign N5366 = ~( N3968 & N4364 );
	assign N6835 = ~( N6566 & N3968 );
	assign N6837 = ~( N6569 & N3968 );
	assign N7871 = ~( N7836 & N3968 );
	assign N7873 = ~( N7839 & N3968 );
	assign N4357 = ~N3968;
	assign OR4_1487_inw1 = ~( N3968 | N5065 );
	assign N4702 = ~( N3810 & N4224 );
	assign N4223 = ~N3810;
	assign N5065 = ( N4357 & N3962 );
	assign N6839 = ~( N6572 & N3962 );
	assign N6841 = ~( N6575 & N3962 );
	assign N7929 = ~( N7900 & N3962 );
	assign N7931 = ~( N7903 & N3962 );
	assign NOR3_1527_inw1 = ~( N3962 | N5117 );
	assign N4364 = ~N3962;
	assign OR4_1526_inw1 = ~( N3962 | N5117 );
	assign N5364 = ~( N3956 & N5108 );
	assign N5106 = ~N3956;
	assign N3908 = ~N3701;
	assign N4701 = ~( N3813 & N4223 );
	assign N4224 = ~N3813;
	assign N5363 = ~( N3948 & N5106 );
	assign N5108 = ~N3948;
	assign N3909 = ~N3702;
	assign N5140 = ~( N3942 & N4855 );
	assign N5110 = ~N3942;
	assign N3914 = ~N3708;
	assign N3975 = ~N3742;
	assign N5371 = ~( N5148 & N5147 );
	assign N5305 = ~( N4008_key & N4405 );
	assign N4521 = ~N4008_key;
	assign N6162 = ( N5606 & N3921 );
	assign N6160 = ~( AND3_1397_inw1 | N3921 );
	assign AND4_1394_inw2 = ~( N3921 & N5264 );
	assign N5137 = ~( N3921 & N4521 );
	assign N6999 = ~( N3921 & N6914 );
	assign N7723 = ~( N7595 & N3921 );
	assign N7782 = ~( N7724 & N3921 );
	assign N4405 = ~N3921;
	assign g16_inw1 = ~( N5579 & N3921 );
	assign N5304 = ~( N3927 & N5113 );
	assign N5115 = ~N3927;
	assign N5303 = ~( N3933 & N5115 );
	assign N5113 = ~N3933;
	assign N5306 = ~( N3732 & N5110 );
	assign N4855 = ~N3732;
	assign N3915 = ~N3709;
	assign N3976 = ~N3743;
	assign AND3_840_inw1 = ~( N3775 & N3771 );
	assign AND3_1003_inw1 = ~( N4188 & N3775 );
	assign N4191 = ~N3775;
	assign N3916 = ~N3710;
	assign N3977 = ~N3744;
	assign AND3_1004_inw1 = ~( N3771 & N4191 );
	assign N4188 = ~N3771;
	assign NOR3_1524_invw = ~( NOR3_1524_inw1 & N6103 );
	assign OR4_1522_inw2 = ~( N6103 | N6133 );
	assign N6100 = ~( AND4_1345_inw1 | AND4_1345_inw2 );
	assign N7080 = ~( N6896 & N6990 );
	assign N6896 = ~( N6553 & N5728 );
	assign N6097 = ~( g12_inw1 | g12_inw2 );
	assign N6138 = ( N5462 & N5452 );
	assign AND3_1374_inw1 = ~( N5462 & N5441 );
	assign AND4_1368_inw1 = ~( N5462 & N5441 );
	assign N7787 = ~( N5462 & N7768 );
	assign N7788 = ~( N5462 & N7770 );
	assign N6651 = ~N5462;
	assign n_305 = ( N5431 & N5462 );
	assign N7076 = ~( N6890 & N6987 );
	assign N6890 = ~( N6536 & N5176 );
	assign N4733 = ~N4109;
	assign AND3_1507_inw1 = ~( N6025 & N4198 );
	assign AND3_1590_inw1 = ~( N4198 & N5315 );
	assign N4524 = ~N4198;
	assign NOR4_1525_invw = ~( NOR4_1525_inw1 & NOR4_1525_inw2 );
	assign g30_inw2 = ~( N6101 | n_316 );
	assign g53_inw2 = ~( N6127 | n_316 );
	assign AND3_1340_inw1 = ~( N5431 & N5424 );
	assign N6099 = ~( AND3_1344_inw1 | N5431 );
	assign AND4_1368_inw2 = ~( N5431 & N5452 );
	assign N6947 = ~( N5431 & N6825 );
	assign N8031 = ~( N5431 & N8020 );
	assign N8032 = ~( N5431 & N8022 );
	assign N6668 = ~N5431;
	assign g2_inw1 = ~( N5441 & N5431 );
	assign g12_inw2 = ~( N5431 & n_307 );
	assign N4736 = ~N4100;
	assign N5155 = ~( N4234 & N4967 );
	assign N4968 = ~N4234;
	assign g10_inw1 = ~( N6095 | N6096 );
	assign N6504 = ~( OR4_1517_inw1 & OR4_1517_inw2 );
	assign N6536 = ~( OR4_1522_inw1 & OR4_1522_inw2 );
	assign AND3_1348_inw1 = ~( N5452 & N5441 );
	assign AND4_1341_inw1 = ~( N5441 & N5424 );
	assign AND4_1345_inw1 = ~( N5452 & N5441 );
	assign AND4_1349_inw2 = ~( N5441 & N5452 );
	assign N6948 = ~( N5441 & N6827 );
	assign N7984 = ~( N5441 & N7966 );
	assign N7985 = ~( N5441 & N7968 );
	assign N6670 = ~N5441;
	assign g8_inw1 = ~( N5441 & N5424 );
	assign n_307 = ( N5452 & N5441 );
	assign g32_inw1 = ~( N5441 & N5452 );
	assign N4735 = ~N4103;
	assign N5154 = ~( N4225 & N4966 );
	assign N4965 = ~N4225;
	assign N6096 = ~( AND4_1341_inw1 | AND4_1341_inw2 );
	assign N7218 = ~( N7080 & N6419 );
	assign N6897 = ~N6419;
	assign N6891 = ( N6419 | N6138 );
	assign N6133 = ~( AND3_1374_inw1 | N5452 );
	assign N6949 = ~( N5452 & N6829 );
	assign N7851 = ~( N5452 & N7832 );
	assign N7852 = ~( N5452 & N7834 );
	assign N6672 = ~N5452;
	assign g8_inw2 = ~( N5452 & n_305 );
	assign N4734 = ~N4106;
	assign N5153 = ~( N4228 & N4965 );
	assign N4966 = ~N4228;
	assign N6084 = ~( AND3_1331_inw1 | N5396 );
	assign N6073 = ~( AND4_1322_inw1 | AND4_1322_inw2 );
	assign N6940 = ~( N6662 & N6816 );
	assign N7212 = ~( N7075 & N7153 );
	assign N6662 = ~( N5407 & N5469 );
	assign N7075 = ~( N6494 & N5469 );
	assign N6089 = ( N5418 & N5407 );
	assign N7176 = ( N5418 & N7023 );
	assign AND3_1332_inw1 = ~( N5418 & N5407 );
	assign AND4_1329_inw1 = ~( N5396 & N5418 );
	assign N7743 = ~( N5418 & N7708 );
	assign N7744 = ~( N5418 & N7710 );
	assign N6079 = ~N5418;
	assign N6939 = ~( N6660 & N6815 );
	assign N7209 = ~( N7073 & N7152 );
	assign N6660 = ~( N5407 & N5087 );
	assign N7073 = ~( N6881 & N5087 );
	assign N4730 = ~N4094;
	assign N5232 = ~( N4240 & N5052 );
	assign N5053 = ~N4240;
	assign g10_inw2 = ~( N6097 | n_306 );
	assign N6946 = ~( N5424 & N6823 );
	assign N7917 = ~( N5424 & N7896 );
	assign N7918 = ~( N5424 & N7898 );
	assign N6666 = ~N5424;
	assign g2_inw2 = ~( N5424 & N6138 );
	assign N4729 = ~N4097;
	assign N5156 = ~( N4231 & N4968 );
	assign N4967 = ~N4231;
	assign N6382 = ~( OR4_1486_inw1 & OR4_1486_inw2 );
	assign AND3_1321_inw1 = ~( N5396 & N5389 );
	assign AND4_1322_inw1 = ~( N5407 & N5389 );
	assign AND4_1329_inw2 = ~( N5407 & N5389 );
	assign N6935 = ~( N5389 & N6807 );
	assign N6936 = ~( N5389 & N6809 );
	assign N7879 = ~( N5389 & N7860 );
	assign N7880 = ~( N5389 & N7862 );
	assign N6653 = ~N5389;
	assign N6066 = ~( N4939 & N5054 );
	assign N5241 = ~N4939;
	assign NOR3_1513_invw = ~( NOR3_1513_inw1 & N6084 );
	assign N6482 = ~( OR4_1512_inw1 & OR4_1512_inw2 );
	assign N6085 = ~( AND3_1332_inw1 | N5396 );
	assign N6937 = ~( N5396 & N6811 );
	assign N6938 = ~( N5396 & N6411 );
	assign N7943 = ~( N5396 & N7924 );
	assign N7944 = ~( N5396 & N7926 );
	assign N6657 = ~N5396;
	assign N4732 = ~N4088;
	assign N6377 = ~( N4243 & N5241 );
	assign N5054 = ~N4243;
	assign OR4_1486_inw2 = ~( N6072 | N6073 );
	assign N6814 = ~( N6494 & N6657 );
	assign N6411 = ~N6494;
	assign N6490 = ~( OR3_1514_inw1 & N6089 );
	assign N7815 = ~( N5407 & N7796 );
	assign N7816 = ~( N5407 & N7798 );
	assign N6661 = ~N5407;
	assign N4731 = ~N4091;
	assign N5233 = ~( N4237 & N5053 );
	assign N5052 = ~N4237;
	assign OR4_1487_inw2 = ~( N5066 | N6074 );
	assign N7087 = ~( N6575 & N5622 );
	assign N6437 = ~N6575;
	assign N6572 = ~( OR3_1528_inw1 & N6147 );
	assign N6147 = ( N5573 & N5562 );
	assign AND3_1383_inw1 = ~( N5573 & N5562 );
	assign AND4_1323_inw1 = ~( N5562 & N4357 );
	assign AND4_1381_inw2 = ~( N5562 & N4357 );
	assign N6689 = ~( N5562 & N5120 );
	assign N6691 = ~( N5562 & N5622 );
	assign N7821 = ~( N5562 & N7806 );
	assign N7822 = ~( N5562 & N7808 );
	assign N6690 = ~N5562;
	assign N5235 = ~( N4144 & N4724 );
	assign N4725 = ~N4144;
	assign N6143 = ~( AND3_1382_inw1 | N4364 );
	assign N6074 = ~( AND4_1323_inw1 | AND4_1323_inw2 );
	assign N6958 = ~( N6691 & N6843 );
	assign N7222 = ~( N7087 & N7159 );
	assign N7181 = ( N5573 & N7049 );
	assign AND4_1381_inw1 = ~( N4364 & N5573 );
	assign N7749 = ~( N5573 & N7718 );
	assign N7750 = ~( N5573 & N7720 );
	assign N6139 = ~N5573;
	assign N6957 = ~( N6689 & N6842 );
	assign N7219 = ~( N7085 & N7158 );
	assign N7085 = ~( N6901 & N5120 );
	assign N5234 = ~( N4147 & N4725 );
	assign N4724 = ~N4147;
	assign g14_inw2 = ~( N6155 | n_308 );
	assign AND3_1390_inw1 = ~( N5264 & N5579 );
	assign AND4_1391_inw1 = ~( N5595 & N5579 );
	assign N6964 = ~( N5579 & N6850 );
	assign N7887 = ~( N5579 & N7874 );
	assign N7923 = ~( N5579 & N7909 );
	assign N6695 = ~N5579;
	assign g4_inw1 = ~( N5595 & N5579 );
	assign g6_inw2 = ~( N5579 & N6194 );
	assign N4728 = ~N4153;
	assign N4975 = ~( N4252 & N4199 );
	assign N4974 = ~N4252;
	assign NOR4_1538_invw = ~( NOR4_1538_inw1 & NOR4_1538_inw2 );
	assign g26_inw2 = ~( N6158 | n_314 );
	assign g51_inw2 = ~( N6184 | n_314 );
	assign N6156 = ~( AND3_1393_inw1 | N5264 );
	assign AND4_1414_inw2 = ~( N5264 & N5606 );
	assign N6965 = ~( N5264 & N6852 );
	assign N8009 = ~( N5264 & N7992 );
	assign N8034 = ~( N5264 & N8026 );
	assign N6434 = ~N5264;
	assign n_303 = ( N5264 & N4405 );
	assign g6_inw1 = ~( N5595 & N5264 );
	assign g16_inw2 = ~( N5264 & n_309 );
	assign N3827 = ~N3456;
	assign g14_inw1 = ~( N6153 | N6154 );
	assign NOR3_1537_invw = ~( NOR3_1537_inw1 & N6160 );
	assign N6584 = ~( OR4_1531_inw1 & OR4_1531_inw2 );
	assign N6606 = ~( OR4_1535_inw1 & OR4_1535_inw2 );
	assign AND3_1397_inw1 = ~( N5606 & N5595 );
	assign AND3_1419_inw1 = ~( N4405 & N5595 );
	assign AND4_1394_inw1 = ~( N5606 & N5595 );
	assign AND4_1398_inw2 = ~( N5595 & N5606 );
	assign AND4_1414_inw1 = ~( N4405 & N5595 );
	assign N6966 = ~( N5595 & N6854 );
	assign N7951 = ~( N5595 & N7938 );
	assign N7987 = ~( N5595 & N7973 );
	assign N6698 = ~N5595;
	assign n_309 = ( N5606 & N5595 );
	assign g28_inw1 = ~( N5595 & N5606 );
	assign N4727 = ~N4156;
	assign N5161 = ~( N4246 & N4973 );
	assign N4972 = ~N4246;
	assign N6154 = ~( AND4_1391_inw1 | AND4_1391_inw2 );
	assign N7229 = ~( N7090 & N6445 );
	assign N6916 = ~N6445;
	assign N6909 = ( N6445 | N6194 );
	assign N6194 = ( N4405 & N5606 );
	assign N6189 = ~( AND3_1419_inw1 | N5606 );
	assign N6699 = ~( N5606 & N5956 );
	assign N7823 = ~( N5606 & N7810 );
	assign N7859 = ~( N5606 & N7845 );
	assign N6700 = ~N5606;
	assign g4_inw2 = ~( N5606 & n_303 );
	assign N4726 = ~N4159;
	assign N5160 = ~( N4249 & N4972 );
	assign N4973 = ~N4249;
	assign N8055 = ~( N8045 & N8033 );
	assign N8056 = ~N8045;
	assign N8013 = ~( OR4_2241_inw1 & OR4_2241_inw2 );
	assign OR4_2241_inw1 = ~( N7988 | N7989 );
	assign OR4_1916_inw1 = ~( N7011 | N7338 );
	assign OR4_1974_inw1 = ~( N7433 | N7434 );
	assign OR4_1976_inw1 = ~( N7339 | N7436 );
	assign OR4_1977_inw1 = ~( N7437 | N7438 );
	assign OR4_1978_inw1 = ~( N7439 | N7440 );
	assign OR4_2088_inw1 = ~( N7666 | N7667 );
	assign OR4_2089_inw1 = ~( N7668 | N7669 );
	assign OR4_2090_inw1 = ~( N7670 | N7671 );
	assign OR4_2091_inw1 = ~( N7672 | N7673 );
	assign OR4_2300_inw1 = ~( N8117 | N8118 );
	assign N7505 = ~( OR4_1974_inw1 & OR4_1974_inw2 );
	assign N7727 = ~( OR4_2088_inw1 & OR4_2088_inw2 );
	assign N7728 = ~( OR4_2089_inw1 & OR4_2089_inw2 );
	assign N7729 = ~( OR4_2090_inw1 & OR4_2090_inw2 );
	assign N7730 = ~( OR4_2091_inw1 & OR4_2091_inw2 );
	assign N7435 = ~( OR4_1916_inw1 & OR4_1916_inw2 );
	assign N7507 = ~( OR4_1976_inw1 & OR4_1976_inw2 );
	assign N7508 = ~( OR4_1977_inw1 & OR4_1977_inw2 );
	assign N7509 = ~( OR4_1978_inw1 & OR4_1978_inw2 );
	assign N8121 = ~( OR4_2300_inw1 & OR4_2300_inw2 );
	assign OR4_1924_inw1 = ~( N7012 | N7340 );
	assign OR4_1979_inw1 = ~( N7441 | N7442 );
	assign OR4_1981_inw1 = ~( N7341 | N7444 );
	assign OR4_1982_inw1 = ~( N7445 | N7446 );
	assign OR4_1983_inw1 = ~( N7447 | N7448 );
	assign OR4_2092_inw1 = ~( N7674 | N7675 );
	assign OR4_2093_inw1 = ~( N7676 | N7677 );
	assign OR4_2094_inw1 = ~( N7678 | N7679 );
	assign OR4_2095_inw1 = ~( N7680 | N7681 );
	assign OR4_2301_inw1 = ~( N8119 | N8120 );
	assign N7510 = ~( OR4_1979_inw1 & OR4_1979_inw2 );
	assign N7731 = ~( OR4_2092_inw1 & OR4_2092_inw2 );
	assign N7732 = ~( OR4_2093_inw1 & OR4_2093_inw2 );
	assign N7733 = ~( OR4_2094_inw1 & OR4_2094_inw2 );
	assign N7734 = ~( OR4_2095_inw1 & OR4_2095_inw2 );
	assign N7443 = ~( OR4_1924_inw1 & OR4_1924_inw2 );
	assign N7512 = ~( OR4_1981_inw1 & OR4_1981_inw2 );
	assign N7513 = ~( OR4_1982_inw1 & OR4_1982_inw2 );
	assign N7514 = ~( OR4_1983_inw1 & OR4_1983_inw2 );
	assign N8122 = ~( OR4_2301_inw1 & OR4_2301_inw2 );
	assign N8057 = ~( N8048 & N8036 );
	assign N8058 = ~N8048;
	assign N8017 = ~( OR4_2242_inw1 & OR4_2242_inw2 );
	assign OR4_2242_inw1 = ~( N7994 | N7995 );
	assign N4273 = ~( OR4_873_inw1 & OR4_873_inw2 );
	assign N4274 = ~( OR4_874_inw1 & OR4_874_inw2 );
	assign N4276 = ~( OR4_876_inw1 & OR4_876_inw2 );
	assign N4277 = ~( OR4_877_inw1 & OR4_877_inw2 );
	assign N7525 = ~( OR4_1992_inw1 & OR4_1992_inw2 );
	assign OR4_1992_inw1 = ~( N4741 | N7114 );
	assign N7449 = ~( OR4_1930_inw1 & OR4_1930_inw2 );
	assign N7736 = ~( OR4_2097_inw1 & OR4_2097_inw2 );
	assign N7737 = ~( OR4_2098_inw1 & OR4_2098_inw2 );
	assign N7738 = ~( OR4_2099_inw1 & OR4_2099_inw2 );
	assign N7739 = ~( OR4_2100_inw1 & OR4_2100_inw2 );
	assign N7515 = ~( OR4_1984_inw1 & OR4_1984_inw2 );
	assign N7516 = ~( OR4_1985_inw1 & OR4_1985_inw2 );
	assign N7517 = ~( OR4_1986_inw1 & OR4_1986_inw2 );
	assign N7518 = ~( OR4_1987_inw1 & OR4_1987_inw2 );
	assign N8123 = ~( OR4_2302_inw1 & OR4_2302_inw2 );
	assign OR4_1930_inw1 = ~( N7013 | N7342 );
	assign OR4_1987_inw1 = ~( N7349 | N7456 );
	assign OR4_1984_inw1 = ~( N7450 | N7451 );
	assign OR4_1985_inw1 = ~( N7452 | N7453 );
	assign OR4_1986_inw1 = ~( N7454 | N7455 );
	assign OR4_2097_inw1 = ~( N7684 | N7685 );
	assign OR4_2098_inw1 = ~( N7686 | N7687 );
	assign OR4_2099_inw1 = ~( N7688 | N7689 );
	assign OR4_2100_inw1 = ~( N7690 | N7691 );
	assign OR4_2302_inw1 = ~( N8113 | N8114 );
	assign OR4_1950_inw1 = ~( N7016 | N7364 );
	assign OR4_1988_inw1 = ~( N7457 | N7458 );
	assign OR4_1989_inw1 = ~( N7459 | N7460 );
	assign OR4_1990_inw1 = ~( N7461 | N7462 );
	assign OR4_1991_inw1 = ~( N7357 | N7463 );
	assign OR4_2096_inw1 = ~( N7682 | N7683 );
	assign OR4_2101_inw1 = ~( N7692 | N7693 );
	assign OR4_2102_inw1 = ~( N7694 | N7695 );
	assign OR4_2103_inw1 = ~( N7696 | N7697 );
	assign OR4_2303_inw1 = ~( N8115 | N8116 );
	assign N7735 = ~( OR4_2096_inw1 & OR4_2096_inw2 );
	assign N7740 = ~( OR4_2101_inw1 & OR4_2101_inw2 );
	assign N7741 = ~( OR4_2102_inw1 & OR4_2102_inw2 );
	assign N7742 = ~( OR4_2103_inw1 & OR4_2103_inw2 );
	assign N7519 = ~( OR4_1988_inw1 & OR4_1988_inw2 );
	assign N7520 = ~( OR4_1989_inw1 & OR4_1989_inw2 );
	assign N7521 = ~( OR4_1990_inw1 & OR4_1990_inw2 );
	assign N7522 = ~( OR4_1991_inw1 & OR4_1991_inw2 );
	assign N8124 = ~( OR4_2303_inw1 & OR4_2303_inw2 );
	assign N7469 = ~( OR4_1950_inw1 & OR4_1950_inw2 );
	assign N8075 = ~( OR4_2278_inw1 & OR4_2278_inw2 );
	assign N8076 = ~( OR4_2279_inw1 & OR4_2279_inw2 );
	assign OR3_1670_inw1 = ~( N4197 | N6718 );
	assign OR3_1837_inw1 = ~( N4956 | N7146 );
	assign OR3_1840_inw1 = ~( N4960 | N7147 );
	assign OR3_1867_inw1 = ~( N4957 | N7187 );
	assign OR3_1868_inw1 = ~( N4958 | N7188 );
	assign OR3_1869_inw1 = ~( N4959 | N7189 );
	assign OR3_1870_inw1 = ~( N4961 | N7196 );
	assign OR3_1871_inw1 = ~( N3998 | N7197 );
	assign OR3_1874_inw1 = ~( N4980 | N7207 );
	assign OR3_1875_inw1 = ~( N4984 | N7208 );
	assign OR3_1998_inw1 = ~( N4981 | N7481 );
	assign OR3_1999_inw1 = ~( N4982 | N7482 );
	assign OR3_2000_inw1 = ~( N4983 | N7483 );
	assign OR3_2001_inw1 = ~( N5165 | N7484 );
	assign OR3_2002_inw1 = ~( N4985 | N7485 );
	assign OR3_2003_inw1 = ~( N4986 | N7486 );
	assign OR3_2004_inw1 = ~( N4547 | N7487 );
	assign OR3_2005_inw1 = ~( N4987 | N7488 );
	assign OR4_2278_inw1 = ~( N7526 | N8071 );
	assign OR4_2279_inw1 = ~( N7636 | N8072 );
	assign N7365 = ~N7190;
	assign N7473 = ~N7270;
	assign N7472 = ~N7276;
	assign N7471 = ~N7282;
	assign N7015 = ~N6866;
	assign N7363 = ~N7198;
	assign N7467 = ~N7288;
	assign N7466 = ~N7294;
	assign N7470 = ~N7304;
	assign N7707 = ~N7531;
	assign N7706 = ~N7537;
	assign N7705 = ~N7543;
	assign N7704 = ~N7549;
	assign N7465 = ~N7310;
	assign N7702 = ~N7555;
	assign N7701 = ~N7561;
	assign N7700 = ~N7567;
	assign N7699 = ~N7573;
	assign N7037 = ~( N6949 & N6830 );
	assign N7245 = ( N7176 | N7040 );
	assign N7236 = ( N7173 | N7125 );
	assign N7239 = ( N7174 | N7126 );
	assign N7242 = ( N7175 | N7127 );
	assign N7173 = ( N7115 & N7023 );
	assign N7174 = ( N7116 & N7023 );
	assign N7175 = ( N6940 & N7023 );
	assign N6828 = ~( N6508 & N6670 );
	assign N6827 = ~N6508;
	assign g33_invw = ~( g33_inw1 & N7034 );
	assign N4278 = N4275;
	assign N6967 = ~( N6699 & N6856 );
	assign N7263 = ( N7181 | N7064 );
	assign N7250 = ( N7178 | N7139 );
	assign N7257 = ( N7179 | N7140 );
	assign N7260 = ( N7180 | N7141 );
	assign N7178 = ( N7130 & N7049 );
	assign N7179 = ( N7131 & N7049 );
	assign N7180 = ( N6958 & N7049 );
	assign N6855 = ~( N6587 & N6698 );
	assign N6854 = ~N6587;
	assign g38_invw = ~( g38_inw1 & N7060 );
	assign N7698 = ( N7624 | N7625 );
	assign N7625 = ( N7489 & N7250 );
	assign N5711 = ~( N5145_key & N5311_key );
	assign N5385 = ~( N5239 & N5059 );
	assign N5707 = ~( N5309_key & N5310_key );
	assign N5703 = ~( N5307_key & N5308_key );
	assign N5331 = ~( N5163 | N4978 );
	assign N5332 = ~( N5164 | N4979 );
	assign N5163 = ~( AND3_1137_inw1 | N4976 );
	assign N5164 = ~( AND3_1138_inw1 | N4976 );
	assign N5236 = ~( N4721 & N5057 );
	assign N4721 = ~( N3911 & N4027 );
	assign N5328 = ~( N5162 & N4975 );
	assign N5060 = ~( AND4_1041_inw1 | AND4_1041_inw2 );
	assign N6475 = ~( AND3_1508_inw1 | N5328 );
	assign N6722 = ~( AND3_1593_inw1 | N6471 );
	assign AND3_1509_inw1 = ~( N6028 & N3987 );
	assign AND3_1592_inw1 = ~( N3987 & N5324 );
	assign N5742 = ~( N5369_key & N5370_key );
	assign AND3_1023_inw1 = ~( N4203 & N4200 );
	assign N5745 = ~( N5367_key & N5368_key );
	assign N5736 = ~( N5365 & N5366_key );
	assign N7044 = ~( N6953 & N6835 );
	assign N7045 = ~( N6954 & N6837 );
	assign N7900 = ~( N7885 & N7871 );
	assign N7903 = ~( N7886 & N7873 );
	assign AND3_1046_inw1 = ~( N4364 & N4357 );
	assign N6953 = ~( N4357 & N6834 );
	assign N6954 = ~( N4357 & N6836 );
	assign N7885 = ~( N4357 & N7870 );
	assign N7886 = ~( N4357 & N7872 );
	assign N6386 = ~( OR4_1487_inw1 & OR4_1487_inw2 );
	assign N5049 = ~( N4701 & N4702 );
	assign N5365 = ~N5065;
	assign N7046 = ~( N6955 & N6839 );
	assign N7047 = ~( N6956 & N6841 );
	assign N7960 = ~( N7945 & N7929 );
	assign N7963 = ~( N7946 & N7931 );
	assign NOR3_1527_invw = ~( NOR3_1527_inw1 & N6143 );
	assign N6144 = ~( AND3_1383_inw1 | N4364 );
	assign N6955 = ~( N4364 & N6838 );
	assign N6956 = ~( N4364 & N6437 );
	assign N7945 = ~( N4364 & N7928 );
	assign N7946 = ~( N4364 & N7930 );
	assign N6566 = ~( OR4_1526_inw1 & OR4_1526_inw2 );
	assign N5739 = ~( N5363_key & N5364_key );
	assign N5700 = ~( N5306_key & N5140_key );
	assign N6024 = ~( N5371 & N5312 );
	assign N6023 = ~N5371;
	assign N5696 = ~( N5137_key & N5305_key );
	assign OR4_1535_inw2 = ~( N6160 | N6189 );
	assign N6157 = ~( AND4_1394_inw1 | AND4_1394_inw2 );
	assign N7090 = ~( N6915 & N6999 );
	assign N7778 = ~( N7751 & N7723 );
	assign N7812 = ~( N7795 & N7782 );
	assign N6915 = ~( N6619 & N4405 );
	assign N7751 = ~( N4405 & N7722 );
	assign N7795 = ~( N4405 & N7781 );
	assign N6155 = ~( g16_inw1 | g16_inw2 );
	assign N5692 = ~( N5303_key & N5304_key );
	assign AND3_1005_inw1 = ~( N4191 & N4188 );
	assign N6553 = ~NOR3_1524_invw;
	assign NOR4_1525_inw2 = ~( N6099 | N6100 );
	assign g30_inw1 = ~( N6099 | N6100 );
	assign g53_inw1 = ~( N6099 | N6100 );
	assign N7217 = ~N7080;
	assign N6127 = ~( AND4_1368_inw1 | AND4_1368_inw2 );
	assign N7800 = ~( N7787 & N7769 );
	assign N7803 = ~( N7788 & N7771 );
	assign N7769 = ~( N7712 & N6651 );
	assign N7771 = ~( N7715 & N6651 );
	assign N7216 = ~( N7076 & N7079 );
	assign N7215 = ~N7076;
	assign AND4_1044_inw1 = ~( N4733 & N4734 );
	assign N6474 = ~( AND3_1507_inw1 | N5319 );
	assign N6719 = ~( AND3_1590_inw1 | N6469 );
	assign AND3_1506_inw1 = ~( N5315 & N4524 );
	assign AND3_1591_inw1 = ~( N4524 & N6025 );
	assign N6556 = ~NOR4_1525_invw;
	assign N6500 = ~( g30_inw1 & g30_inw2 );
	assign N6539 = ~( g53_inw1 & g53_inw2 );
	assign N7031 = ~( N6947 & N6826 );
	assign N8037 = ~( N8031 & N8021 );
	assign N8038 = ~( N8032 & N8023 );
	assign N6826 = ~( N6504 & N6668 );
	assign N8021 = ~( N7998 & N6668 );
	assign N8023 = ~( N8001 & N6668 );
	assign N6117 = ~( g2_inw1 | g2_inw2 );
	assign AND4_1044_inw2 = ~( N4735 & N4736 );
	assign N5319 = ~( N5155 & N5156 );
	assign N6397 = ~( g10_inw1 & g10_inw2 );
	assign N6825 = ~N6504;
	assign N6889 = ~N6536;
	assign N7034 = ~( N6948 & N6828 );
	assign N7998 = ~( N7984 & N7967 );
	assign N8001 = ~( N7985 & N7969 );
	assign N7967 = ~( N7932 & N6670 );
	assign N7969 = ~( N7935 & N6670 );
	assign N6091 = ~( g8_inw1 | g8_inw2 );
	assign N5315 = ~( N5153 & N5154 );
	assign N7412 = ~( N7321 & N7218 );
	assign N7321 = ~( N6897 & N7217 );
	assign N7320 = ~( N6891 & N7215 );
	assign N7079 = ~N6891;
	assign N7864 = ~( N7851 & N7833 );
	assign N7867 = ~( N7852 & N7835 );
	assign N7833 = ~( N7800 & N6672 );
	assign N7835 = ~( N7803 & N6672 );
	assign OR4_1512_inw2 = ~( N6084 | N6085 );
	assign N7408 = ~( N7212 & N6809 );
	assign N7407 = ~N7212;
	assign N6881 = ( N6411 | N6089 );
	assign N6080 = ~( AND4_1329_inw1 | AND4_1329_inw2 );
	assign N7762 = ~( N7743 & N7709 );
	assign N7765 = ~( N7744 & N7711 );
	assign N7709 = ~( N7579 & N6079 );
	assign N7711 = ~( N7582 & N6079 );
	assign N7022 = ~N6939;
	assign N7406 = ~( N7209 & N6807 );
	assign N7405 = ~N7209;
	assign AND4_1043_inw1 = ~( N4729 & N4730 );
	assign N5377 = ~( N5232 & N5233 );
	assign N7028 = ~( N6946 & N6824 );
	assign N7932 = ~( N7917 & N7897 );
	assign N7935 = ~( N7918 & N7899 );
	assign N6824 = ~( N6500 & N6666 );
	assign N7897 = ~( N7864 & N6666 );
	assign N7899 = ~( N7867 & N6666 );
	assign N6924 = ( N6382 | N6801 );
	assign N7018 = ~( N6935 & N6808 );
	assign N7019 = ~( N6936 & N6810 );
	assign N7890 = ~( N7879 & N7861 );
	assign N7893 = ~( N7880 & N7863 );
	assign N6808 = ~( N6482 & N6653 );
	assign N6810 = ~( N6486 & N6653 );
	assign N7861 = ~( N7826 & N6653 );
	assign N7863 = ~( N7829 & N6653 );
	assign N6634 = ~( N6377 & N6066 );
	assign N5388 = ~( AND3_1237_inw1 | N5241 );
	assign N6486 = ~NOR3_1513_invw;
	assign N7492 = ~( N6482 & N7405 );
	assign N6807 = ~N6482;
	assign N7020 = ~( N6937 & N6812 );
	assign N7021 = ~( N6938 & N6814 );
	assign N7954 = ~( N7943 & N7925 );
	assign N7957 = ~( N7944 & N7927 );
	assign N6812 = ~( N6490 & N6657 );
	assign N7925 = ~( N7890 & N6657 );
	assign N7927 = ~( N7893 & N6657 );
	assign AND4_1043_inw2 = ~( N4731 & N4732 );
	assign N6811 = ~N6490;
	assign N7826 = ~( N7815 & N7797 );
	assign N7829 = ~( N7816 & N7799 );
	assign N7797 = ~( N7762 & N6661 );
	assign N7799 = ~( N7765 & N6661 );
	assign N6901 = ( N6437 | N6147 );
	assign N6838 = ~N6572;
	assign N6140 = ~( AND4_1381_inw1 | AND4_1381_inw2 );
	assign N7836 = ~( N7821 & N7807 );
	assign N7839 = ~( N7822 & N7809 );
	assign N7807 = ~( N7772 & N6690 );
	assign N7809 = ~( N7775 & N6690 );
	assign N5382 = ~( N5234 & N5235 );
	assign AND4_1041_inw1 = ~( N4724 & N4725 );
	assign OR4_1526_inw2 = ~( N6143 | N6144 );
	assign N7418 = ~( N7222 & N6836 );
	assign N7417 = ~N7222;
	assign N7772 = ~( N7749 & N7719 );
	assign N7775 = ~( N7750 & N7721 );
	assign N7719 = ~( N7589 & N6139 );
	assign N7721 = ~( N7592 & N6139 );
	assign N7048 = ~N6957;
	assign N7416 = ~( N7219 & N6834 );
	assign N7415 = ~N7219;
	assign N6427 = ~( g14_inw1 & g14_inw2 );
	assign N7054 = ~( N6964 & N6851 );
	assign N7906 = ~( N7887 & N7875 );
	assign N7940 = ~( N7923 & N7910 );
	assign N6851 = ~( N6580 & N6695 );
	assign N7875 = ~( N7842 & N6695 );
	assign N7910 = ~( N7876 & N6695 );
	assign N6149 = ~( g4_inw1 | g4_inw2 );
	assign N6175 = ~( g6_inw1 | g6_inw2 );
	assign AND4_1042_inw2 = ~( N3827 & N4728 );
	assign N6622 = ~NOR4_1538_invw;
	assign N6580 = ~( g26_inw1 & g26_inw2 );
	assign N6609 = ~( g51_inw1 & g51_inw2 );
	assign NOR4_1538_inw2 = ~( N6156 | N6157 );
	assign g26_inw1 = ~( N6156 | N6157 );
	assign g51_inw1 = ~( N6156 | N6157 );
	assign N6184 = ~( AND4_1414_inw1 | AND4_1414_inw2 );
	assign N7057 = ~( N6965 & N6853 );
	assign N8025 = ~( N8009 & N7993 );
	assign N8039 = ~( N8034 & N8027 );
	assign N6853 = ~( N6584 & N6434 );
	assign N7993 = ~( N7970 & N6434 );
	assign N8027 = ~( N8004 & N6434 );
	assign N6619 = ~NOR3_1537_invw;
	assign N6852 = ~N6584;
	assign N7160 = ~( N6606 & N7088 );
	assign N6912 = ~N6606;
	assign N7060 = ~( N6966 & N6855 );
	assign N7970 = ~( N7951 & N7939 );
	assign N8004 = ~( N7987 & N7974 );
	assign N7939 = ~( N7906 & N6698 );
	assign N7974 = ~( N7940 & N6698 );
	assign AND4_1042_inw1 = ~( N4726 & N4727 );
	assign N5324 = ~( N5160 & N5161 );
	assign N7421 = ~( N7328 & N7229 );
	assign N7328 = ~( N6916 & N7228 );
	assign N7089 = ~( N6909 & N6912 );
	assign N7088 = ~N6909;
	assign N7842 = ~( N7823 & N7811 );
	assign N7876 = ~( N7859 & N7846 );
	assign N7811 = ~( N7778 & N6700 );
	assign N7846 = ~( N7812 & N6700 );
	assign N8061 = ~( N8055 & N8059 );
	assign N8059 = ~( N8013 & N8056 );
	assign N8033 = ~N8013;
	assign N8064 = ~( N8057 & N8060 );
	assign N8060 = ~( N8017 & N8058 );
	assign N8036 = ~N8017;
	assign n_320 = ~( N7245 | N7242 );
	assign n_321 = ~( N7239 | N7236 );
	assign n_318 = ~g33_invw;
	assign n_325 = ~( N7263 | N7260 );
	assign N7432 = ~N7250;
	assign n_322 = ~N7257;
	assign n_323 = ~g38_invw;
	assign N6714 = ~( AND3_1586_inw1_key | N5711_key );
	assign N6715 = ~( AND3_1587_inw1_key | N5711_key );
	assign N6710 = ~N5711_key;
	assign N6477 = ~( N5385 & N6234 );
	assign N6044 = ~N5385;
	assign AND3_1586_inw1 = ~( N5707_key & N5703_key );
	assign AND3_1668_inw1 = ~( N6203 & N5707_key );
	assign N6206 = ~N5707_key;
	assign AND3_1669_inw1 = ~( N5703_key & N6206 );
	assign N6203 = ~N5703_key;
	assign N5756 = ~( N5332 & N5331 );
	assign N6378 = ~( N5236 & N6068 );
	assign N5755 = ~N5236;
	assign N6476 = ~( AND3_1509_inw1 | N5328 );
	assign N6471 = ~N5328;
	assign AND3_1175_inw1 = ~( N5060 & N5061 );
	assign N6874 = ~( N6721 | N6475 );
	assign N6875 = ~( N6722 | N6476 );
	assign N6721 = ~( AND3_1592_inw1 | N6471 );
	assign N6633 = ~( N5742_key & N6376 );
	assign N6375 = ~N5742_key;
	assign N6632 = ~( N5745_key & N6375 );
	assign N6376 = ~N5745_key;
	assign N6631 = ~( N5736_key & N6374 );
	assign N6373 = ~N5736_key;
	assign N7130 = ~N7045;
	assign N7928 = ~N7900;
	assign N7930 = ~N7903;
	assign N6925 = ( N6386 | N6802 );
	assign N6221 = ~( N5049 & N6023 );
	assign N5312 = ~N5049;
	assign N7131 = ~N7047;
	assign AND3_2234_inw1 = ~( N7960 & N6427 );
	assign AND3_2236_inw1 = ~( N7960 & N7182 );
	assign AND3_2233_inw1 = ~( N7963 & N6857 );
	assign AND3_2235_inw1 = ~( N7963 & N7065 );
	assign N6569 = ~NOR3_1527_invw;
	assign N7498 = ~( N6566 & N7415 );
	assign N6834 = ~N6566;
	assign N6630 = ~( N5739_key & N6373 );
	assign N6374 = ~N5739_key;
	assign N6712 = ~( AND3_1584_inw1_key | N5700_key );
	assign N6713 = ~( AND3_1585_inw1_key | N5700_key );
	assign N6708 = ~N5700_key;
	assign N6716 = ~( N6221 & N6024 );
	assign AND3_1584_inw1 = ~( N5696_key & N5692_key );
	assign AND3_1666_inw1 = ~( N6197 & N5696_key );
	assign N6200 = ~N5696_key;
	assign N7228 = ~N7090;
	assign N7810 = ~N7778;
	assign N7845 = ~N7812;
	assign AND3_1667_inw1 = ~( N5692_key & N6200 );
	assign N6197 = ~N5692_key;
	assign N6895 = ~N6553;
	assign N7832 = ~N7800;
	assign N7834 = ~N7803;
	assign N7409 = ~( N7320 & N7216 );
	assign N5063 = ~( AND4_1044_inw1 | AND4_1044_inw2 );
	assign N6873 = ~( N6720 | N6474 );
	assign N6872 = ~( N6719 | N6473 );
	assign N6473 = ~( AND3_1506_inw1 | N5319 );
	assign N6720 = ~( AND3_1591_inw1 | N6469 );
	assign N7658 = ~( N6556 & N7587 );
	assign N6900 = ~N6556;
	assign N6823 = ~N6500;
	assign N7657 = ~( N6539 & N7585 );
	assign N6894 = ~N6539;
	assign n_319 = ~( N7031 | N7028 );
	assign N8040 = ~N8038;
	assign N6641 = ( N6080 & N6117 );
	assign N6675 = ~N6117;
	assign N6469 = ~N5319;
	assign N6801 = ( N6080 & N6397 );
	assign AND3_2228_inw1 = ~( N7954 & N6397 );
	assign N6831 = ~N6397;
	assign N8020 = ~N7998;
	assign N8022 = ~N8001;
	assign N6648 = ( N6080 & N6091 );
	assign N6025 = ~N5315;
	assign N7588 = ~( N7412 & N6900 );
	assign N7587 = ~N7412;
	assign N7896 = ~N7864;
	assign N7898 = ~N7867;
	assign N7582 = ~( N7493 & N7408 );
	assign N7493 = ~( N6486 & N7407 );
	assign N7072 = ~N6881;
	assign N7796 = ~N7762;
	assign N7798 = ~N7765;
	assign N7579 = ~( N7492 & N7406 );
	assign N5062 = ~( AND4_1043_inw1 | AND4_1043_inw2 );
	assign N7002 = ~( N5377 & N6922 );
	assign N6067 = ~N5377;
	assign N7966 = ~N7932;
	assign N7968 = ~N7935;
	assign N6926 = N6924;
	assign N7115 = ~N7019;
	assign N7924 = ~N7890;
	assign N7926 = ~N7893;
	assign N6923 = ~( N6634 & N6067 );
	assign N6922 = ~N6634;
	assign N6809 = ~N6486;
	assign N7116 = ~N7021;
	assign AND3_2230_inw1 = ~( N7954 & N7177 );
	assign AND3_2227_inw1 = ~( N7957 & N6831 );
	assign AND3_2229_inw1 = ~( N7957 & N7041 );
	assign N7860 = ~N7826;
	assign N7862 = ~N7829;
	assign N7084 = ~N6901;
	assign N6643 = ( N6140 & N6149 );
	assign N6646 = ( N6140 & N6175 );
	assign N6802 = ( N6427 & N6140 );
	assign N7870 = ~N7836;
	assign N7872 = ~N7839;
	assign N6069 = ~( N5382 & N5755 );
	assign N6068 = ~N5382;
	assign N7592 = ~( N7499 & N7418 );
	assign N7499 = ~( N6569 & N7417 );
	assign N7806 = ~N7772;
	assign N7808 = ~N7775;
	assign N7589 = ~( N7498 & N7416 );
	assign N6857 = ~N6427;
	assign n_324 = ~( N7057 | N7054 );
	assign N7938 = ~N7906;
	assign N7973 = ~N7940;
	assign N6703 = ~N6175;
	assign N5061 = ~( AND4_1042_inw1 | AND4_1042_inw2 );
	assign N7665 = ~( N6622 & N7598 );
	assign N6919 = ~N6622;
	assign N6850 = ~N6580;
	assign N7500 = ~( N6609 & N7419 );
	assign N6913 = ~N6609;
	assign N8042 = ~N8039;
	assign N6914 = ~N6619;
	assign N7225 = ~( N7089 & N7160 );
	assign N7992 = ~N7970;
	assign N8026 = ~N8004;
	assign N6028 = ~N5324;
	assign N7599 = ~( N7421 & N6919 );
	assign N7598 = ~N7421;
	assign N7874 = ~N7842;
	assign N7909 = ~N7876;
	assign N8073 = ~N8061;
	assign N8074 = ~N8064;
	assign g37_inw2 = ~( n_320 & n_321 );
	assign g37_inw1 = ~( n_318 & n_319 );
	assign g43_inw2 = ~( n_325 & n_326 );
	assign n_326 = ( n_322 & N7432 );
	assign g43_inw1 = ~( n_323 & n_324 );
	assign N6975 = ~( N6862_key | N6714_key );
	assign N6976 = ~( N6863_key | N6715_key );
	assign N6862 = ~( AND3_1668_inw1_key | N6710 );
	assign N6863 = ~( AND3_1669_inw1_key | N6710 );
	assign N6877 = ~( N6477 & N6235 );
	assign N6235 = ~( N5756 & N6044 );
	assign AND3_1587_inw1 = ~( N6206 & N6203 );
	assign N6234 = ~N5756;
	assign N6637 = ~( N6069 & N6378 );
	assign N7006 = ~( N6875 & N6874 );
	assign N6795 = ~( N6632_key & N6633_key );
	assign N6792 = ~( N6630_key & N6631_key );
	assign N6927 = N6925;
	assign N6836 = ~N6569;
	assign N6973 = ~( N6860_key | N6712_key );
	assign N6974 = ~( N6861_key | N6713_key );
	assign N6860 = ~( AND3_1666_inw1_key | N6708 );
	assign N6861 = ~( AND3_1667_inw1_key | N6708 );
	assign g44_invw = ~( g44_inw1_key & N6716 );
	assign AND3_1585_inw1 = ~( N6200 & N6197 );
	assign N7586 = ~( N7409 & N6894 );
	assign N7585 = ~N7409;
	assign AND3_1237_inw1 = ~( N5062 & N5063 );
	assign N7003 = ~( N6873 & N6872 );
	assign N7715 = ~( N7658 & N7588 );
	assign N7712 = ~( N7657 & N7586 );
	assign N7041 = ( N6831 & N6675 );
	assign N7710 = ~N7582;
	assign N7708 = ~N7579;
	assign N7101 = ~( N7002 & N6923 );
	assign N7720 = ~N7592;
	assign N7718 = ~N7589;
	assign N7065 = ( N6857 & N6703 );
	assign N7724 = ~( N7665 & N7599 );
	assign N7595 = ~( N7500 & N7420 );
	assign N7420 = ~( N7225 & N6913 );
	assign N7419 = ~N7225;
	assign N7503 = ~( g37_inw1 | g37_inw2 );
	assign N7504 = ~( g43_inw1 | g43_inw2 );
	assign N7097 = ~( N6976_key & N6975_key );
	assign n_327 = ~N6877;
	assign N7206 = ~( N6637 & N7150 );
	assign N6876 = ~N6637;
	assign N7151 = ~( N7006 & N6876 );
	assign N7150 = ~N7006;
	assign N7269 = ~( N6795_key & N7185 );
	assign N6978 = ~N6795_key;
	assign N7268 = ~( N6792_key & N7183 );
	assign N6977 = ~N6792_key;
	assign N7094 = ~( N6974_key & N6973_key );
	assign n_328 = ~g44_invw;
	assign N7300 = ~( N7003 & N7205 );
	assign N7149 = ~N7003;
	assign N7770 = ~N7715;
	assign N7768 = ~N7712;
	assign N7177 = ~N7041;
	assign N7204 = ~( N7101 & N7149 );
	assign N7205 = ~N7101;
	assign N7182 = ~N7065;
	assign N7781 = ~N7724;
	assign N7722 = ~N7595;
	assign N7186 = ~( N7097_key & N6978 );
	assign N7185 = ~N7097_key;
	assign N7301 = ~( N7206 & N7151 );
	assign N7476 = ~( N7269_key & N7186_key );
	assign N7474 = ~( N7268_key & N7184_key );
	assign N7184 = ~( N7094_key & N6977 );
	assign N7183 = ~N7094_key;
	assign N7402 = ~( N7204_key & N7300_key );
	assign N7468 = ~N7301_key;
	assign g44_inw1 = ~( N7474_key | N7476_key );
	assign N7529 = ~N7402_key;
	assign g44_inw1_key = ~( g44_inw1 ^ key_0 );
	assign N7402_key = ~( N7402 ^ key_1 );
	assign N7184_key = ~( N7184 ^ key_2 );
	assign N7474_key = ~( N7474 ^ key_3 );
	assign N7476_key = ~( N7476 ^ key_4 );
	assign N7301_key = ~( N7301 ^ key_5 );
	assign N7186_key = ~( N7186 ^ key_6 );
	assign N7204_key = ~( N7204 ^ key_7 );
	assign N7300_key = ~( N7300 ^ key_8 );
	assign N7094_key = ~( N7094 ^ key_9 );
	assign N7268_key = ~( N7268 ^ key_10 );
	assign N7269_key = ~( N7269 ^ key_11 );
	assign N372_key = ~( N372 ^ key_12 );
	assign N2954_key = ~( N2954 ^ key_13 );
	assign N3723_key = ~( N3723 ^ key_14 );
	assign N4008_key = ~( N4008 ^ key_15 );
	assign N5366_key = ~( N5366 ^ key_16 );
	assign N5364_key = ~( N5364 ^ key_17 );
	assign N5363_key = ~( N5363 ^ key_18 );
	assign N5140_key = ~( N5140 ^ key_19 );
	assign N5305_key = ~( N5305 ^ key_20 );
	assign N5137_key = ~( N5137 ^ key_21 );
	assign N5304_key = ~( N5304 ^ key_22 );
	assign N5303_key = ~( N5303 ^ key_23 );
	assign N5306_key = ~( N5306 ^ key_24 );
	assign N5736_key = ~( N5736 ^ key_25 );
	assign N5739_key = ~( N5739 ^ key_26 );
	assign N5700_key = ~( N5700 ^ key_27 );
	assign N5696_key = ~( N5696 ^ key_28 );
	assign N5692_key = ~( N5692 ^ key_29 );
	assign N6631_key = ~( N6631 ^ key_30 );
	assign N6630_key = ~( N6630 ^ key_31 );
	assign N6712_key = ~( N6712 ^ key_32 );
	assign N6713_key = ~( N6713 ^ key_33 );
	assign AND3_1584_inw1_key = ~( AND3_1584_inw1 ^ key_34 );
	assign AND3_1666_inw1_key = ~( AND3_1666_inw1 ^ key_35 );
	assign AND3_1667_inw1_key = ~( AND3_1667_inw1 ^ key_36 );
	assign N6792_key = ~( N6792 ^ key_37 );
	assign N6973_key = ~( N6973 ^ key_38 );
	assign N6974_key = ~( N6974 ^ key_39 );
	assign N6860_key = ~( N6860 ^ key_40 );
	assign N6861_key = ~( N6861 ^ key_41 );
	assign AND3_1585_inw1_key = ~( AND3_1585_inw1 ^ key_42 );
	assign N292_key = ~( N292 ^ key_43 );
	assign N3680_key = ~( N3680 ^ key_44 );
	assign N2867_key = ~( N2867 ^ key_45 );
	assign N4011_key = ~( N4011 ^ key_46 );
	assign N5145_key = ~( N5145 ^ key_47 );
	assign N5310_key = ~( N5310 ^ key_48 );
	assign N5309_key = ~( N5309 ^ key_49 );
	assign N5308_key = ~( N5308 ^ key_50 );
	assign N5307_key = ~( N5307 ^ key_51 );
	assign N5370_key = ~( N5370 ^ key_52 );
	assign N5369_key = ~( N5369 ^ key_53 );
	assign N5368_key = ~( N5368 ^ key_54 );
	assign N5367_key = ~( N5367 ^ key_55 );
	assign N5311_key = ~( N5311 ^ key_56 );
	assign N5711_key = ~( N5711 ^ key_57 );
	assign N5707_key = ~( N5707 ^ key_58 );
	assign N5703_key = ~( N5703 ^ key_59 );
	assign N5742_key = ~( N5742 ^ key_60 );
	assign N5745_key = ~( N5745 ^ key_61 );
	assign N6714_key = ~( N6714 ^ key_62 );
	assign N6715_key = ~( N6715 ^ key_63 );
	assign AND3_1586_inw1_key = ~( AND3_1586_inw1 ^ key_64 );
	assign AND3_1668_inw1_key = ~( AND3_1668_inw1 ^ key_65 );
	assign AND3_1669_inw1_key = ~( AND3_1669_inw1 ^ key_66 );
	assign N6633_key = ~( N6633 ^ key_67 );
	assign N6632_key = ~( N6632 ^ key_68 );
	assign N6975_key = ~( N6975 ^ key_69 );
	assign N6976_key = ~( N6976 ^ key_70 );
	assign N6862_key = ~( N6862 ^ key_71 );
	assign N6863_key = ~( N6863 ^ key_72 );
	assign AND3_1587_inw1_key = ~( AND3_1587_inw1 ^ key_73 );
	assign N6795_key = ~( N6795 ^ key_74 );
	assign N7097_key = ~( N7097 ^ key_75 );
	assign N566_key = ~( N566 ^ key_76 );
	assign N3027_key = ~( N3027 ^ key_77 );
	assign N3023_key = ~( N3023 ^ key_78 );
	assign N3028_key = ~( N3028 ^ key_79 );
	assign N3024_key = ~( N3024 ^ key_80 );
	assign N3029_key = ~( N3029 ^ key_81 );
	assign N3025_key = ~( N3025 ^ key_82 );
	assign N3030_key = ~( N3030 ^ key_83 );
	assign N3026_key = ~( N3026 ^ key_84 );
	assign N2938_key = ~( N2938 ^ key_85 );
	assign N2939_key = ~( N2939 ^ key_86 );
	assign N2940_key = ~( N2940 ^ key_87 );
	assign N2941_key = ~( N2941 ^ key_88 );
	assign AND3_377_inw1_key = ~( AND3_377_inw1 ^ key_89 );
	assign AND3_378_inw1_key = ~( AND3_378_inw1 ^ key_90 );
	assign AND3_379_inw1_key = ~( AND3_379_inw1 ^ key_91 );
	assign AND3_380_inw1_key = ~( AND3_380_inw1 ^ key_92 );
	assign AND3_444_inw1_key = ~( AND3_444_inw1 ^ key_93 );
	assign AND3_445_inw1_key = ~( AND3_445_inw1 ^ key_94 );
	assign AND3_446_inw1_key = ~( AND3_446_inw1 ^ key_95 );
	assign AND3_447_inw1_key = ~( AND3_447_inw1 ^ key_96 );
	assign AND3_524_inw1_key = ~( AND3_524_inw1 ^ key_97 );
	assign AND3_525_inw1_key = ~( AND3_525_inw1 ^ key_98 );
	assign AND3_526_inw1_key = ~( AND3_526_inw1 ^ key_99 );
	assign AND3_527_inw1_key = ~( AND3_527_inw1 ^ key_100 );
	assign AND3_547_inw1_key = ~( AND3_547_inw1 ^ key_101 );
	assign AND3_548_inw1_key = ~( AND3_548_inw1 ^ key_102 );
	assign AND3_549_inw1_key = ~( AND3_549_inw1 ^ key_103 );
	assign AND3_550_inw1_key = ~( AND3_550_inw1 ^ key_104 );
	assign N3463_key = ~( N3463 ^ key_105 );
	assign N3464_key = ~( N3464 ^ key_106 );
	assign N3465_key = ~( N3465 ^ key_107 );
	assign N3466_key = ~( N3466 ^ key_108 );
	assign N3508_key = ~( N3508 ^ key_109 );
	assign N3509_key = ~( N3509 ^ key_110 );
	assign N3510_key = ~( N3510 ^ key_111 );
	assign N3511_key = ~( N3511 ^ key_112 );
	assign N2934_key = ~( N2934 ^ key_113 );
	assign N2935_key = ~( N2935 ^ key_114 );
	assign N2936_key = ~( N2936 ^ key_115 );
	assign N2937_key = ~( N2937 ^ key_116 );
	assign N4608_key = ~( N4608 ^ key_117 );
	assign N3722_key = ~( N3722 ^ key_118 );
	assign N3719_key = ~( N3719 ^ key_119 );
	assign N3720_key = ~( N3720 ^ key_120 );
	assign N3721_key = ~( N3721 ^ key_121 );
	assign N3769_key = ~( N3769 ^ key_122 );
	assign N3770_key = ~( N3770 ^ key_123 );
endmodule
