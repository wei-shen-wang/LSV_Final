module c432(N1, N102, N105, N108, N11, N112, N115, N14, N17, N21, N24, N27, N30, N34, N37, N4, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N8, N82, N86, N89, N92, N95, N99, key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, N223, N329, N370, N421, N430, N431, N432);
	input N1, N102, N105, N108, N11, N112, N115, N14, N17, N21, N24, N27, N30, N34, N37, N4, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N8, N82, N86, N89, N92, N95, N99;
	input key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12;
	output N223, N329, N370, N421, N430, N431, N432;
	wire N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N242, N118, N154, NAND4_138_inw1, N119, N334, N157, N246, N122, N371, N158, N159, NAND4_139_inw2, N123, N336, N183, N250, N126, N372, N184, N162, NAND4_140_inw2, N127, N338, N185, N254, N130, N373, N186, N165, NAND4_141_inw2, N131, N340, N187, N255, N134, N374, N188, N168, NAND4_142_inw2, N135, N342, N189, N256, N138, N375, N190, N171, NAND4_143_inw2, N139, N344, N191, N257, N142, N376, N192, N174, NAND4_144_inw2, N143, N345, N193, N258, N146, N377, N194, N177, NAND4_145_inw2, N147, N346, N195, N259, N150, N378, N196, N180, NAND4_146_inw2, N151, N347, N197, N379, N198, N224, g1_inw1, NAND4_138_invw, NAND4_138_inw2, N260, NAND4_139_inw1, N263, N227, NAND4_139_invw, N264, NAND4_140_inw1, N288, N230, n_44, NAND4_140_invw, N267, NAND4_141_inw1, N289, N233, n_45, NAND4_141_invw, N270, NAND4_142_inw1, N290, N236, NAND4_142_invw, N273, NAND4_143_inw1, N291, N239, n_46, NAND4_143_invw, N276, NAND4_144_inw1, N292, N243, NAND4_144_invw, N279, NAND4_145_inw1, N293, N247, n_47, NAND4_145_invw, N282, NAND4_146_inw1, N294, N251, NAND4_146_invw, N285, N295, N380, N330, g6_inw1, N300, N381, N331, N301, g5_inw1, N386, N332, n_48, N302, N393, N333, n_49, N303, N399, N335, N304, g5_inw2, N404, N337, n_50, N305, N407, N339, N306, N411, N341, n_51, N307, N414, N343, N308, N415, N348, NAND4_158_inw1, NAND4_159_inw1, NAND4_160_inw1, n_56, N349, N199, N422, NAND4_155_inw1, NAND4_157_inw1, N350, g10_inw1, NAND3_156_inw1, N417, n_57, N351, NAND4_155_inw2, NAND4_158_inw2, N352, N418, n_58, N353, g10_inw2, NAND4_157_inw2, N419, N354, N420, n_59, N355, N356, N421, g11_inw1, NAND4_158_invw, NAND4_159_invw, NAND4_160_invw, g20_inw1, N223, NAND4_155_invw, NAND4_157_invw, n_52, N296, NAND3_156_invw, n_53, g20_inw2, n_54, n_55, N430, N431, N432, N416, N425, N429, g15_inw1, N329, N428, g15_inw2, NAND4_159_inw2, NAND4_160_inw2, N357, N370;
	wire N357_key, NAND4_160_inw2_key, N14_key, N27_key, N40_key, N53_key, N66_key, N79_key, N92_key, N105_key, N115_key, N158_key, N184_key;
	wire key_0, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12;
	assign N242 = ~( N1 & N223 );
	assign N118 = ~N1;
	assign N154 = ~( N118 & N4 );
	assign NAND4_138_inw1 = ~( N4 & N242 );
	assign N119 = ~N4;
	assign N334 = ~( N8 & N329 );
	assign N157 = ~( N8 | N119 );
	assign N246 = ~( N223 & N11 );
	assign N122 = ~N11;
	assign N371 = ~( N14_key & N370 );
	assign N158 = ~( N14_key | N119 );
	assign N159 = ~( N122 & N17 );
	assign NAND4_139_inw2 = ~( N372 & N17 );
	assign N123 = ~N17;
	assign N336 = ~( N329 & N21 );
	assign N183 = ~( N21 | N123 );
	assign N250 = ~( N223 & N24 );
	assign N126 = ~N24;
	assign N372 = ~( N370 & N27_key );
	assign N184 = ~( N27_key | N123 );
	assign N162 = ~( N126 & N30 );
	assign NAND4_140_inw2 = ~( N373 & N30 );
	assign N127 = ~N30;
	assign N338 = ~( N329 & N34 );
	assign N185 = ~( N34 | N127 );
	assign N254 = ~( N223 & N37 );
	assign N130 = ~N37;
	assign N373 = ~( N370 & N40_key );
	assign N186 = ~( N40_key | N127 );
	assign N165 = ~( N130 & N43 );
	assign NAND4_141_inw2 = ~( N374 & N43 );
	assign N131 = ~N43;
	assign N340 = ~( N329 & N47 );
	assign N187 = ~( N47 | N131 );
	assign N255 = ~( N223 & N50 );
	assign N134 = ~N50;
	assign N374 = ~( N370 & N53_key );
	assign N188 = ~( N53_key | N131 );
	assign N168 = ~( N134 & N56 );
	assign NAND4_142_inw2 = ~( N375 & N56 );
	assign N135 = ~N56;
	assign N342 = ~( N329 & N60 );
	assign N189 = ~( N60 | N135 );
	assign N256 = ~( N223 & N63 );
	assign N138 = ~N63;
	assign N375 = ~( N370 & N66_key );
	assign N190 = ~( N66_key | N135 );
	assign N171 = ~( N138 & N69 );
	assign NAND4_143_inw2 = ~( N376 & N69 );
	assign N139 = ~N69;
	assign N344 = ~( N329 & N73 );
	assign N191 = ~( N73 | N139 );
	assign N257 = ~( N223 & N76 );
	assign N142 = ~N76;
	assign N376 = ~( N370 & N79_key );
	assign N192 = ~( N79_key | N139 );
	assign N174 = ~( N142 & N82 );
	assign NAND4_144_inw2 = ~( N377 & N82 );
	assign N143 = ~N82;
	assign N345 = ~( N329 & N86 );
	assign N193 = ~( N86 | N143 );
	assign N258 = ~( N223 & N89 );
	assign N146 = ~N89;
	assign N377 = ~( N370 & N92_key );
	assign N194 = ~( N92_key | N143 );
	assign N177 = ~( N146 & N95 );
	assign NAND4_145_inw2 = ~( N378 & N95 );
	assign N147 = ~N95;
	assign N346 = ~( N329 & N99 );
	assign N195 = ~( N99 | N147 );
	assign N259 = ~( N223 & N102 );
	assign N150 = ~N102;
	assign N378 = ~( N370 & N105_key );
	assign N196 = ~( N105_key | N147 );
	assign N180 = ~( N150 & N108 );
	assign NAND4_146_inw2 = ~( N379 & N108 );
	assign N151 = ~N108;
	assign N347 = ~( N329 & N112 );
	assign N197 = ~( N112 | N151 );
	assign N379 = ~( N370 & N115_key );
	assign N198 = ~( N115_key | N151 );
	assign N224 = ( N223 ^ N154 );
	assign g1_inw1 = ~( N154 & N159 );
	assign NAND4_138_invw = ~( NAND4_138_inw1 | NAND4_138_inw2 );
	assign NAND4_138_inw2 = ~( N334 & N371 );
	assign N260 = ~( N224 & N157 );
	assign NAND4_139_inw1 = ~( N246 & N336 );
	assign N263 = ~( N224 & N158_key );
	assign N227 = ( N223 ^ N159 );
	assign NAND4_139_invw = ~( NAND4_139_inw1 | NAND4_139_inw2 );
	assign N264 = ~( N227 & N183 );
	assign NAND4_140_inw1 = ~( N250 & N338 );
	assign N288 = ~( N227 & N184_key );
	assign N230 = ( N223 ^ N162 );
	assign n_44 = ~( g1_inw1 | N162 );
	assign NAND4_140_invw = ~( NAND4_140_inw1 | NAND4_140_inw2 );
	assign N267 = ~( N230 & N185 );
	assign NAND4_141_inw1 = ~( N254 & N340 );
	assign N289 = ~( N230 & N186 );
	assign N233 = ( N223 ^ N165 );
	assign n_45 = ( N165 & N168 );
	assign NAND4_141_invw = ~( NAND4_141_inw1 | NAND4_141_inw2 );
	assign N270 = ~( N233 & N187 );
	assign NAND4_142_inw1 = ~( N255 & N342 );
	assign N290 = ~( N233 & N188 );
	assign N236 = ( N223 ^ N168 );
	assign NAND4_142_invw = ~( NAND4_142_inw1 | NAND4_142_inw2 );
	assign N273 = ~( N236 & N189 );
	assign NAND4_143_inw1 = ~( N256 & N344 );
	assign N291 = ~( N236 & N190 );
	assign N239 = ( N223 ^ N171 );
	assign n_46 = ( N171 & N174 );
	assign NAND4_143_invw = ~( NAND4_143_inw1 | NAND4_143_inw2 );
	assign N276 = ~( N239 & N191 );
	assign NAND4_144_inw1 = ~( N257 & N345 );
	assign N292 = ~( N239 & N192 );
	assign N243 = ( N223 ^ N174 );
	assign NAND4_144_invw = ~( NAND4_144_inw1 | NAND4_144_inw2 );
	assign N279 = ~( N243 & N193 );
	assign NAND4_145_inw1 = ~( N258 & N346 );
	assign N293 = ~( N243 & N194 );
	assign N247 = ( N223 ^ N177 );
	assign n_47 = ( N177 & N180 );
	assign NAND4_145_invw = ~( NAND4_145_inw1 | NAND4_145_inw2 );
	assign N282 = ~( N247 & N195 );
	assign NAND4_146_inw1 = ~( N259 & N347 );
	assign N294 = ~( N247 & N196 );
	assign N251 = ( N223 ^ N180 );
	assign NAND4_146_invw = ~( NAND4_146_inw1 | NAND4_146_inw2 );
	assign N285 = ~( N251 & N197 );
	assign N295 = ~( N251 & N198 );
	assign N380 = ~NAND4_138_invw;
	assign N330 = ( N329 ^ N260 );
	assign g6_inw1 = ~( N260 & N264 );
	assign N300 = ~N263;
	assign N381 = ~NAND4_139_invw;
	assign N331 = ( N329 ^ N264 );
	assign N301 = ~N288;
	assign g5_inw1 = ~( n_44 & n_45 );
	assign N386 = ~NAND4_140_invw;
	assign N332 = ( N329 ^ N267 );
	assign n_48 = ~( g6_inw1 | N267 );
	assign N302 = ~N289;
	assign N393 = ~NAND4_141_invw;
	assign N333 = ( N329 ^ N270 );
	assign n_49 = ( N270 & N273 );
	assign N303 = ~N290;
	assign N399 = ~NAND4_142_invw;
	assign N335 = ( N329 ^ N273 );
	assign N304 = ~N291;
	assign g5_inw2 = ~( n_46 & n_47 );
	assign N404 = ~NAND4_143_invw;
	assign N337 = ( N329 ^ N276 );
	assign n_50 = ( N276 & N279 );
	assign N305 = ~N292;
	assign N407 = ~NAND4_144_invw;
	assign N339 = ( N329 ^ N279 );
	assign N306 = ~N293;
	assign N411 = ~NAND4_145_invw;
	assign N341 = ( N329 ^ N282 );
	assign n_51 = ( N282 & N285 );
	assign N307 = ~N294;
	assign N414 = ~NAND4_146_invw;
	assign N343 = ( N329 ^ N285 );
	assign N308 = ~N295;
	assign N415 = ~N380;
	assign N348 = ~( N330 & N300 );
	assign NAND4_158_inw1 = ~( N381 & N386 );
	assign NAND4_159_inw1 = ~( N381 & N386 );
	assign NAND4_160_inw1 = ~( N381 & N422 );
	assign n_56 = ( N381 & N386 );
	assign N349 = ~( N331 & N301 );
	assign N199 = ~( g5_inw1 | g5_inw2 );
	assign N422 = ~( N386 & N417 );
	assign NAND4_155_inw1 = ~( N386 & N393 );
	assign NAND4_157_inw1 = ~( N386 & N393 );
	assign N350 = ~( N332 & N302 );
	assign g10_inw1 = ~( n_48 & n_49 );
	assign NAND3_156_inw1 = ~( N399 & N393 );
	assign N417 = ~N393;
	assign n_57 = ( N393 & N399 );
	assign N351 = ~( N333 & N303 );
	assign NAND4_155_inw2 = ~( N418 & N399 );
	assign NAND4_158_inw2 = ~( N422 & N399 );
	assign N352 = ~( N335 & N304 );
	assign N418 = ~N404;
	assign n_58 = ( N404 & N407 );
	assign N353 = ~( N337 & N305 );
	assign g10_inw2 = ~( n_50 & n_51 );
	assign NAND4_157_inw2 = ~( N407 & N420 );
	assign N419 = ~N407;
	assign N354 = ~( N339 & N306 );
	assign N420 = ~N411;
	assign n_59 = ( N411 & N414 );
	assign N355 = ~( N341 & N307 );
	assign N356 = ~( N343 & N308 );
	assign N421 = ~( N415 | N416 );
	assign g11_inw1 = ~( N348 & N349 );
	assign NAND4_158_invw = ~( NAND4_158_inw1 | NAND4_158_inw2 );
	assign NAND4_159_invw = ~( NAND4_159_inw1 | NAND4_159_inw2 );
	assign NAND4_160_invw = ~( NAND4_160_inw1 | NAND4_160_inw2_key );
	assign g20_inw1 = ~( n_56 & n_57 );
	assign N223 = ~N199;
	assign NAND4_155_invw = ~( NAND4_155_inw1 | NAND4_155_inw2 );
	assign NAND4_157_invw = ~( NAND4_157_inw1 | NAND4_157_inw2 );
	assign n_52 = ~( g11_inw1 | N350 );
	assign N296 = ~( g10_inw1 | g10_inw2 );
	assign NAND3_156_invw = ~( NAND3_156_inw1 | N419 );
	assign n_53 = ( N351 & N352 );
	assign g20_inw2 = ~( n_58 & n_59 );
	assign n_54 = ( N353 & N354 );
	assign n_55 = ( N355 & N356 );
	assign N430 = ~NAND4_158_invw;
	assign N431 = ~NAND4_159_invw;
	assign N432 = ~NAND4_160_invw;
	assign N416 = ~( g20_inw1 | g20_inw2 );
	assign N425 = ~NAND4_155_invw;
	assign N429 = ~NAND4_157_invw;
	assign g15_inw1 = ~( n_52 & n_53 );
	assign N329 = ~N296;
	assign N428 = ~NAND3_156_invw;
	assign g15_inw2 = ~( n_54 & n_55 );
	assign NAND4_159_inw2 = ~( N425 & N428 );
	assign NAND4_160_inw2 = ~( N425 & N429 );
	assign N357 = ~( g15_inw1 | g15_inw2 );
	assign N370 = ~N357_key;
	assign N357_key = ~( N357 ^ key_0 );
	assign NAND4_160_inw2_key = ~( NAND4_160_inw2 ^ key_1 );
	assign N14_key = ~( N14 ^ key_2 );
	assign N27_key = ~( N27 ^ key_3 );
	assign N40_key = ~( N40 ^ key_4 );
	assign N53_key = ~( N53 ^ key_5 );
	assign N66_key = ~( N66 ^ key_6 );
	assign N79_key = ~( N79 ^ key_7 );
	assign N92_key = ~( N92 ^ key_8 );
	assign N105_key = ~( N105 ^ key_9 );
	assign N115_key = ~( N115 ^ key_10 );
	assign N158_key = ~( N158 ^ key_11 );
	assign N184_key = ~( N184 ^ key_12 );
endmodule
