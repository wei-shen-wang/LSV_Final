module c7552(N1, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N12, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N15, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N18, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N23, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241_I, N242, N245, N248, N251, N254, N257, N26, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N29, N293, N296, N299, N303, N307, N310, N313, N316, N319, N32, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N35, N352, N355, N358, N361, N364, N367, N38, N382, N41, N44, N47, N5, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N9, N94, N97, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N1110, N1111, N1112, N1113, N1114, N11333, N11334, N11340, N11342, N1489, N1490, N1781, N241_O, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945);
	input N1, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N12, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N15, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N18, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N23, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241_I, N242, N245, N248, N251, N254, N257, N26, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N29, N293, N296, N299, N303, N307, N310, N313, N316, N319, N32, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N35, N352, N355, N358, N361, N364, N367, N38, N382, N41, N44, N47, N5, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N9, N94, N97;
	output N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N1110, N1111, N1112, N1113, N1114, N11333, N11334, N11340, N11342, N1489, N1490, N1781, N241_O, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945;
	wire N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N1490, N889, N388, N387, N1781, N585, N628, N582, N1782, N1793, N1794, N1795, N1796, N1797, N1798, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2337, N2338, N2339, N2340, N2341, N2374, N2375, N2376, N2377, N2378, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N3005, N3006, N3007, N3008, N3009, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N695, N2674, N2680, N1930, N1929, N1928, N2012, N2011, N1167, N1537, N1649, N1966, N2107, N2268, N2355, N2653, N1708, N1822, N1927, N1926, N2010, N2013, N2424, N2425, N2426, N2427, N467, N2396, N2399, N2403, N2404, N2405, N2434, N2433, N2429, N2014, N2418, N2367, N2423, N2420, N2422, N2421, N2397, N2398, N2402, N2401, N2400, N2428, N2430, N2431, N2432, N2435, N2361, N2363, AND4_2717_inw1, N9407, n_333, N2324, N2323, N2303, N2299, N945, N4467, N674, N2436, N2437, N2360, N2362, N2359, N2358, N2321, N2322, N2325, N2302, N2301, N2300, N469, N2281, N2279, N2277, N2280, N2278, AND4_21_inw1, AND4_42_inw1, AND4_11_inw1, AND4_41_inw1, AND4_41_inw2, AND4_11_inw2, AND4_42_inw2, AND4_21_inw2, N1110, N2364, N641, N478, N642, N643, N4471, N644, N482, N4469, N651, N484, N4465, N660, N486, N4463, N666, N489, N688, N672, N492, N700, N673, N2365, N705, N501, N706, N707, N4523, N708, N505, N4519, N715, N507, N4517, N721, N509, N4515, N727, N511, N4513, N599, N513, N4521, N734, N515, N4511, N742, N517, N4509, N604, N519, N4507, N609, N535, N758, N537, N759, N539, N5958, N762, N541, N5956, N768, N543, N5954, N774, N545, N5952, N780, N547, N5950, N786, N549, N5948, N794, N551, N5946, N800, N553, N5944, N806, N556, N812, N813, N6076, N814, N559, N6074, N821, N561, N6072, N827, N563, N6070, N833, N565, N6068, N839, N567, N6066, N845, N569, N6064, N853, N571, N6062, N859, N573, N6060, N865, N9288, N9767, N11316, AND3_2476_inw1, AND3_2853_inw1, AND3_2863_inw1, N11224, N11225, AND4_2475_inw1, AND4_2851_inw1, AND4_2861_inw1, N9773, N9893, N1115, n_318, n_353, N1028, N1029, N241_O, N1109, N881, N2441, N2446, N2450, N2454, N2458, N2462, N2466, N2470, N2474, N2478, N2482, N2488, N2496, N2502, N2508, N2619, N2626, N2632, N2638, N2644, N2766, N2769, N2772, N2775, N4490, N4496, N5322, N3073, g43_inw1, N1114, N1111, N2239, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2793, N2538, N2542, N2546, N2550, N2778, N2554, N2561, N2567, N2573, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2781, N2654, N2658, N2662, N2666, N2670, N2787, N2784, N2796, N2729, N2733, N2737, N2741, N2745, N2749, N2753, N2757, N2761, N2790, N2604, N2607, N2611, N2615, N2688, N2692, N2696, N2700, N2704, N3247, N3251, N3255, N3259, N3263, N3267, N3273, N3281, N3287, N3293, N3789, N3299, N3303, N3307, N3311, N3783, N3315, N3322, N3328, N3334, N3786, N3340, N3343, N3349, N3355, N3384, N3390, N3398, N3404, N3410, N3891, N3416, N3420, N3424, N3428, N3432, N3436, N3440, N3444, N3448, N3888, N3885, N3454, N3458, N3462, N3466, N3470, N3474, N3478, N3482, N2366, N3381, N4769, N5960, N7744, N6217, N4575, N6690, N4768, n_350, N3507, OR3_922_inw1, N2866, N4488, N6712, N2537, N4193, N3379, N2257, N2523, N2650, N2988, N4487, N6711, N2117, N2108, N2111, N2172, N2357, N9790, N9817, g34_inw2, N5654, N3101, N5169, N528, N578, N494, N575, N1112, N5683, N3114, N5171, N3515, N5670, N3107, N5170, N5640, N3097, N5168, N5632, N3096, N5167, N957, N1821, N5856, N3202, N5204, N3628, N5837, N3195, N5202, N5821, N3189, N5201, N5807, N3185, N5200, N5799, N3184, N5199, N5850, N3178, N5203, N3625, N5789, N3173, N5198, N5778, N3169, N5197, N5771, N3168, N5196, N6957, N4570, N6547, N6946, N4566, N6546, N6936, N4563, N6545, N6929, N4562, N6544, N6923, N4555, N6543, N4844, N6912, N4549, N6542, N6901, N4545, N6541, N6894, N4544, N6540, N7180, N4687, N6629, N5030, N7170, N4682, N6628, N7159, N4678, N6627, N7149, N4675, N6626, N7142, N4674, N6625, N7136, N4667, N6624, N4940, N7125, N4661, N6623, N7114, N4657, N6622, N7107, N4656, N6621, N9635, g87_inw2, N9925, N11323, N9287, N10043, N10061, OR4_3452_inw2, N9286, N10041, N10059, N9932, N10025, N11308, N11222, N11223, N9740, g5_inw2, g75_inw2, N1222, N2171, N1113, N3080, N3373, N5185, N5320, N4498, N5186, N5318, N4497, g40_inw2, N3371, N5187, N5316, N4500, N3370, N5188, N5314, N4499, N3365, N5289, N5433, N4618, N3364, N5297, N5584, N4626, N5287, N5585, N4616, g44_inw2, N3362, N5285, N5586, N4614, N3361, N5283, N5587, N4612, N5193, N4505, N5474, N4522, N5475, N4512, N5476, N4510, N5477, N4508, N4472, N5180, N4470, N5181, N4468, N5182, N4466, N5183, N4464, N4327, N3551, N4326, N3552, N4334, N3569, N4333, N3570, N5736, N5747, N6059, N5179, N5184, N5323, N7106, N5429, N3453, N4751, N5299, N4628, g62_inw1, N3368, N5295, N5430, N4624, N5293, N5431, N4622, g59_inw2, N3366, N5291, N5432, N4620, N5189, N3167, N4502, N4501, N5190, N4504, N5191, N4503, N5192, N4506, N5363, N3380, N4694, N4651, n_338, N5321, N5364, N4649, N5319, N5365, N4647, N5317, N5366, N4645, N5315, N5367, N4643, N4411, N3782, N4412, N3781, N5451, N3486, N4776, N5300, N4627, n_346, N5296, N5452, N4623, N5294, N5453, N4621, N5292, N5454, N4619, N5290, N5455, N4617, N5298, N5602, N4625, N5288, N5603, N4615, N5286, N5604, N4613, N5284, N5605, N4611, N5425, N3452, N4746, N4745, N4766, N5426, N6687, N4748, N5427, N6686, N4747, g67_inw2, N4762, N6668, N6685, N4749, N4637, N6597, N6661, N4636, N4635, N5571, N6604, N4642, N5572, N6596, N4633, g53_inw2, N4632, N5573, N6595, N4631, N4630, N5574, N6594, N4629, N4760, N6136, N6683, N6135, N4759, N6688, N6741, N6163, N6681, N6742, N6153, g56_inw2, N4757, N6679, N6743, N6151, N4756, N6677, N6744, N6149, N6648, N5953, N6733, N5951, N6734, N5949, N6735, N5947, N6736, N5945, N6658, N4743, N6122, N6605, N6040, g66_inw1, N4640, N6602, N6659, N6036, N6600, N6660, N6034, g63_inw2, N4638, N6125, N6598, N6032, N6639, N4699, N6091, N6077, N6640, N6075, N6641, N6073, N6642, N6071, N6644, N4700, N6097, N6096, N6645, N5959, N6646, N5957, N6647, N5955, N6643, N6069, N6729, N6067, N6730, N6065, N6731, N6063, N6732, N6061, N6706, N4783, N6186, N6606, N6039, n_348, N6603, N6707, N6035, N6601, N6708, N6033, N6599, N6709, N6031, N6030, N6710, N6029, N6038, N6755, N6037, N6028, N6756, N6027, N6026, N6757, N6025, N6024, N6758, N6023, N5456, N4782, N5457, N4781, N6161, N6702, N6160, N6159, N6703, N6158, N6157, N6704, N6156, N6684, N6705, N6154, N6689, N6751, N6162, N6682, N6752, N6152, N6680, N6753, N6150, N6678, N6754, N6148, N6164, N6165, g70_inw1, N6967, N6968, N8357, N8356, AND4_2115_inw2, N9863, N8717, g29_inw1, N8326, N10086, N7552, N7377, g70_inw2, N5165, N6194, N9065, N3126, N4303, N5178, N7444, N3955, N10451, N5324, n_331, N3122, N3953, N10271, N10272, N3954, N10731, N9955, N9956, N3135, N3375, N5177, N7441, N6192, OR4_2905_inw2, N10054, N10053, N9734, N6777, AND3_1756_inw1, AND3_1763_inw1, AND3_1764_inw1, AND4_1753_inw1, AND4_1757_inw1, AND4_1758_inw1, AND4_2965_inw2, N10644, N11141, N11142, N8250, n_320, g11_inw1, g77_inw1, g95_inw1, N6770, N6767, NOR3_2032_inw1, OR4_2030_inw1, OR4_3029_inw1, N886, N882, N883, N887, N885, N884, N6783, N10281, AND3_2966_inw1, AND4_2965_inw1, N10565, N10737, N10738, N8247, n_321, N6782, N6778, AND4_1757_inw2, N9435, N6195, N10428, g9_inw1, N9432, N4795, N6779, N10280, AND4_1758_inw2, N10645, N10909, N10910, N8251, g11_inw2, AND4_1753_inw2, N7613, OR3_3030_inw1, AND3_1752_inw1, N6771, N10643, N11242, N11243, N8249, g9_inw2, g95_inw2, N6766, NOR4_2033_inw1, n_362, N10642, N11023, N11024, N8248, g77_inw2, n_319, N6866, N10290, AND3_1816_inw1, AND3_2972_inw1, AND4_1810_inw1, AND4_2971_inw1, N10552, N10746, N10747, N8242, n_322, N6864, N6860, AND4_1809_inw2, N9445, N6203, N10415, g25_inw1, N9442, N4813, AND3_1815_inw1, N6861, N10289, AND4_1809_inw1, AND4_1810_inw2, AND4_2971_inw2, N10640, N10915, N10916, N8246, g13_inw2, n_328, g91_inw1, N6859, AND3_1808_inw1, AND4_1805_inw2, N7659, OR3_3026_inw1, AND4_1805_inw1, N10639, N11143, N11144, N8245, g13_inw1, g79_inw1, N6852, N6849, NOR3_2040_inw1, OR4_2038_inw1, OR4_3025_inw1, AND3_1804_inw1, N6853, N10638, N11244, N11245, N8244, g25_inw2, g91_inw2, N6848, NOR4_2041_inw1, n_360, N10637, N11027, N11028, N8243, g79_inw2, n_325, N6865, N10710, AND3_1798_inw1, AND4_1792_inw1, N10609, N10610, N6761, N6844, AND3_1797_inw1, AND4_1795_inw2, N8888, N9847, N5943, N8887, N9846, N4543, AND4_1795_inw1, N8322, N8324, N10845, N10846, N8323, N6839, N6837, N8208, OR3_2044_inw1, AND3_1794_inw1, N6840, N6841, AND4_1792_inw2, N9273, N9274, N11077, N11078, N8294, N6836, NOR3_2037_inw1, OR4_2036_inw1, N9271, N9272, N10969, N10970, N8315, OR4_2019_inw1, N9318, AND3_2117_inw1, N9315, AND4_2115_inw1, AND4_2475_inw2, AND4_2488_inw2, N10035, N10981, N11031, N9252, g17_inw2, n_330, g87_inw1, N8355, AND3_2114_inw1, AND4_2111_inw2, N8931, OR3_2646_inw1, AND3_2489_inw1, AND4_2111_inw1, AND4_2488_inw1, N10034, N11210, N11250, N9251, g17_inw1, g83_inw1, N8352, N8349, NOR3_2424_inw1, OR4_2645_inw1, OR4_2667_inw1, AND3_2110_inw1, N8353, N10033, N11282, N11295, N9250, n_324, g29_inw2, N8348, NOR4_2425_inw1, n_358, N10032, N11095, N11145, N9249, g83_inw2, n_327, N8346, N10269, AND3_2103_inw1, AND4_2097_inw1, N10748, N10749, N8253, N8345, AND3_2102_inw1, AND4_2100_inw2, N9570, N10085, N6969, N9569, N10084, N5966, AND4_2097_inw2, AND4_2100_inw1, N9297, N9299, N10917, N10918, N9298, N8340, N8338, N9111, OR3_2420_inw1, AND3_2099_inw1, N8341, N8342, N9764, N9765, N11137, N11138, N9294, N8337, NOR3_2419_inw1, OR4_2418_inw1, N9762, N9763, N11029, N11030, N9290, OR4_2371_inw1, N8518, N10597, AND3_2217_inw1, AND3_3108_inw1, AND4_2211_inw1, AND4_3107_inw1, N10764, N10862, N10863, N9244, n_323, N8456, N8455, AND4_2177_inw2, N9876, N7573, N10668, g27_inw1, N9873, N6235, AND3_2179_inw1, N8513, N10596, AND4_2177_inw1, AND4_2211_inw2, AND4_3107_inw2, N10835, N10986, N10987, N9248, g15_inw2, n_329, g99_inw1, N8454, AND3_2176_inw1, AND4_2173_inw2, N9005, OR3_3136_inw1, AND4_2173_inw1, N10834, N11211, N11212, N9247, g15_inw1, g81_inw1, N8451, N8448, NOR3_2440_inw1, OR4_2438_inw1, OR4_3135_inw1, AND3_2172_inw1, N8452, N10833, N11284, N11285, N9246, g27_inw2, g99_inw2, N8447, NOR4_2441_inw1, n_364, N10832, N11098, N11099, N9245, g81_inw2, n_326, N8442, N10867, AND3_2164_inw1, AND4_2158_inw1, N10753, N10754, N8252, N8441, AND3_2163_inw1, AND4_2161_inw2, N9601, N10094, N7187, N9600, N10093, N6078, AND4_2158_inw2, AND4_2161_inw1, N9359, N9361, N10922, N10923, N9360, N8436, N8434, N9173, OR3_2430_inw1, AND3_2160_inw1, N8437, N8438, N9797, N9798, N11139, N11140, N9356, N8433, NOR3_2429_inw1, OR4_2428_inw1, N9795, N9796, N11034, N11035, N9352, OR4_2382_inw1, N9904, N9903, N9285, N10105, N10106, N10107, N10108, N10130, N10124, N11336, N11337, N9632, N10119, N10148, N11252, OR4_2645_inw2, OR4_2892_inw2, OR4_2906_inw2, N10133, N10131, OR4_3452_inw1, N10015, N10022, N1489, AND4_1887_inw2, N5751, N6056, N6052, N7104, N7103, N5755, N6047, n_334, N6041, n_342, N6003, N6145, AND4_1869_inw2, N6021, N6252, N6000, N7061, N7060, N5996, N6249, OR4_2027_inw1, N5991, N5766, N6199, N6196, N5740, N5744, N4803, N4806, AND3_2075_inw1, AND3_2353_inw1, N6797, AND3_2077_inw1, AND3_2355_inw1, N6803, n_339, g36_inw2, N6137, N6022, N7067, AND4_1873_inw2, N6018, N6141, N6014, N7065, N7064, N6009, N5758, N5762, N6079, g43_inw2, N6083, N6087, N4997, N6166, g62_inw2, N6170, N6174, N6266, N6263, N6127, AND4_2240_inw2, N6131, N7373, N7369, N8552, N8551, N7331, N7364, n_343, N7080, N7322, AND4_2151_inw2, N6246, N7098, N7077, N8410, N8409, N6243, N7073, OR4_2378_inw1, N7068, n_344, N7358, AND4_2236_inw2, N7376, N7577, N7355, N8546, N8545, N7351, N7574, OR4_2392_inw1, N7346, N7213, N7569, N7566, N7314, N7099, N8418, AND4_2155_inw2, N7095, N7318, N7091, N8416, N8415, N7086, N7194, N7198, N7202, N7205, N7209, N7563, N7560, N7394, g66_inw2, N7398, N7402, N7591, N7588, N6177, N7387, N7391, N7585, N7582, N8554, NOR3_2424_invw, OR4_2667_inw2, N8354, N9979, N9691, N8351, N10857, N10919, N9741, N10192, N9976, n_341, N10549, N10631, N9429, N10551, N10705, N8610, N4784, n_316, N9064, N5469, N10730, N8609, N10628, N5631, g32_inw2, N8262, N8269, N8818, N4473, N10357, N10360, N10212, N10213, N10839, N10070, N10073, N10588, N9836, N9838, N8421, N8960, N4653, N5735, N8608, N8607, N10140, N10233, N10139, g32_inw1, N6768, N6772, N6773, N10279, N10717, N11168, N11171, N10571, N11115, N11117, N6784, N6762, N10278, g7_inw1, NOR3_2032_invw, N8114, N10422, AND3_3130_inw1, N9068, N10641, N10789, N10792, N10466, N10672, N10674, OR4_2030_inw2, OR4_3029_inw2, N9646, N9073, N10573, N10572, N6769, N9642, N9067, N10425, N10718, N10928, N10931, N10873, N10875, N9960, N9074, NOR4_2033_inw2, g93_inw1, g103_inw1, N10716, N11260, N11261, N10569, N11214, N11216, NOR4_2033_invw, g93_inw2, g103_inw2, N10715, N11044, N11047, N10567, N10989, N10991, g7_inw2, N9089, N6855, N10288, N10632, N10800, N10803, N10456, N10682, N10684, NOR3_2040_invw, OR4_2038_inw2, OR4_3025_inw2, N6854, N9667, N9094, N10564, N10563, N6851, N9663, N9088, N10412, N10714, N10938, N10941, N10883, N10885, N6881, N10287, N6850, N9970, N9095, N10713, N11174, N11177, N10562, N11119, N11121, N6845, g19_inw1, N8166, N10409, NOR4_2041_inw2, g89_inw1, g101_inw1, N10712, N11262, N11263, N10560, N11218, N11220, NOR4_2041_invw, g89_inw2, g101_inw2, N10711, N11050, N11053, N10558, N10999, N11001, g19_inw2, N9079, N8204, N10763, N6833, N10675, N10678, N10556, N10516, N10518, N6838, N9243, N9964, N9662, N9275, N9961, N9660, N10876, N10879, N10797, N10799, OR4_2019_inw2, N8886, N7650, NOR3_2037_invw, OR4_2036_inw2, N9540, N9556, N11100, N11103, N8884, N11041, N11043, N8146, N9539, N9555, N10992, N10995, N8880, N8882, N10935, N10937, N7649, N9682, N9314, N10112, N11008, N11062, N10954, N11007, N9280, N8350, N10196, N9692, N10111, N11233, N11272, N9902, N11184, N11232, N9307, g23_inw1, N9629, N9679, NOR4_2425_inw2, g85_inw1, g107_inw1, N10110, N11292, N11307, N9900, N11265, N11291, NOR4_2425_invw, g85_inw2, g107_inw2, N10109, N11124, N11180, N9898, N11066, N11123, g23_inw2, N9671, N9107, N10353, N8333, N10806, N10809, N10686, N10688, N8339, N9742, N10189, N9974, N9766, N10186, N9972, N10944, N10947, N10887, N10889, OR4_2371_inw2, N9568, N8924, NOR3_2419_invw, OR4_2418_inw2, N9895, N9924, N11156, N11159, N9566, N11107, N11109, N9099, N9894, N9923, N11056, N11059, N9562, N9564, N11003, N11005, N8898, N9717, N8507, N10595, N10827, N10899, N10902, N10720, N10824, N10826, NOR3_2440_invw, OR4_2438_inw2, OR4_3135_inw2, N8453, N10003, N9722, N10776, N10775, N8450, N9999, N9716, N10665, N10871, N11015, N11018, N10962, N10964, N8444, N10594, N8449, N10206, N9723, N10870, N11236, N11239, N10774, N11186, N11188, N8497, g21_inw1, N9203, N10662, NOR4_2441_inw2, g97_inw1, g105_inw1, N10869, N11293, N11294, N10772, N11268, N11270, NOR4_2441_invw, g97_inw2, g105_inw2, N10868, N11127, N11130, N10770, N11074, N11076, g21_inw2, N9707, N9169, N10908, N8430, N10817, N10820, N10768, N10695, N10697, N8435, N9739, N10200, N9998, N9799, N10197, N9996, N10955, N10958, N10896, N10898, OR4_2382_inw2, N9599, N8996, NOR3_2429_invw, OR4_2428_inw2, N9891, N9946, N11162, N11165, N9597, N11111, N11113, N9161, N9890, N9945, N11067, N11070, N9593, N9595, N11012, N11014, N8963, N10350, N10351, N10352, N10381, N10266, N10267, N10268, N10292, N11341, N11339, N9901, N11280, N11154, N11155, N10283, N10291, N10455, N11283, N10116, N10141, N10301, N10230, g3_inw1, g73_inw1, N7105, AND3_2354_inw1, N6806, n_337, AND4_1887_inw1, g46_inw1, g36_inw1, N8282, N8283, N8276, g40_inw1, g46_inw2, g52_inw2, AND4_1873_inw1, g39_inw1, g59_inw1, N8539, N8540, N8537, N7062, AND4_1866_inw1, N8216, N7557, AND4_1869_inw1, OR4_2027_inw2, AND4_1866_inw2, g44_inw1, N8217, N7556, N7825, N8284, N8285, N8278, N8144, N7478, N8145, N7477, AND3_2352_inw1, N6800, N8280, N8281, N8274, N10036, N5769, N10037, N5770, N8862, AND3_2076_inw1, N8864, AND3_2078_inw1, N7852, AND3_2231_inw1, AND3_2391_inw1, N7334, n_335, N7066, n_336, AND3_2390_inw1, N7337, g52_inw1, AND3_2079_inw1, AND3_2357_inw1, N6809, AND3_2356_inw1, N6812, AND3_2191_inw1, AND3_2385_inw1, N7188, AND3_2384_inw1, N7191, N8483, N8484, N8469, N10062, N6102, AND3_2251_inw1, AND3_2395_inw1, N7378, AND3_2394_inw1, N7381, N8578, N8579, N8564, N8232, N7581, N8233, N7580, AND3_2531_inw1, AND3_2636_inw1, N7325, N8553, AND3_2635_inw1, N7328, n_349, AND4_2240_inw1, g50_inw1, g58_inw1, N9398, N9399, N9394, g67_inw1, g55_inw2, AND4_2155_inw1, g48_inw2, g63_inw1, N9396, N9397, N9392, N8411, N8218, N7559, AND4_2148_inw1, AND4_2151_inw1, OR4_2378_inw2, N8219, N7558, AND4_2148_inw2, g53_inw1, N8950, g58_inw2, g50_inw2, N8547, AND4_2233_inw1, N9159, N8734, AND4_2236_inw1, OR4_2392_inw2, AND4_2233_inw2, g56_inw1, N9160, N8733, N9029, N9371, N9372, N9365, N9181, N8756, N9182, N8755, AND3_2529_inw1, AND3_2634_inw1, N8519, n_340, N8417, n_347, AND3_2633_inw1, N8522, g48_inw1, g55_inw1, AND3_2515_inw1, AND3_2628_inw1, N8457, AND3_2627_inw1, N8460, N9369, N9370, N9363, AND3_2517_inw1, AND3_2630_inw1, N8463, AND3_2629_inw1, N8466, N9179, N8754, N9180, N8753, AND3_2547_inw1, AND3_2643_inw1, N8558, AND3_2642_inw1, N8561, N9421, N9422, N9415, N9234, N8815, N9235, N8814, AND3_2545_inw1, AND3_2641_inw1, N7384, AND3_2640_inw1, N8555, N9419, N9420, N9413, N9236, N8817, N9237, N8816, N9146, N10195, N10892, N10950, N10816, N10891, N10333, N10332, N10759, N10706, N9837, N6191, g3_inw2, g73_inw2, N9426, N10837, N10546, N10102, N9736, N10020, AND4_2835_inw2, N9732, N10013, AND4_2828_inw2, AND3_3101_inw1, AND3_3132_inw1, AND3_3100_inw1, AND3_3131_inw1, N10840, N10241, N10242, N9526, N10016, AND4_2831_inw2, N10587, N10234, N10295, N11213, N11215, N10282, N10270, N8254, N7609, N8131, N9066, N10568, N10647, N10076, N9645, N10872, N10874, N9959, N9958, N9957, N10570, N10988, N10990, N10173, N10077, N10419, N8117, N11278, N11277, N8134, N11114, N11116, N10082, N9666, N10882, N10884, N8183, N9969, N9968, N9967, N10561, N10998, N11000, N8307, N10183, N10083, N11217, N11219, N8298, N8288, N7655, N9087, N10559, N10406, N8169, N11279, N8186, N11118, N11120, N9659, N8883, N8874, N10796, N10798, N10709, N10179, N10178, N9541, N10177, N10176, N10934, N10936, N8156, N10554, N9738, AND3_3403_inw1, AND3_3405_inw1, AND3_3402_inw1, AND3_3404_inw1, N10247, N8879, N10553, N9737, N11040, N11042, N9265, N10441, N9977, N11065, N11122, N9754, N10334, N10259, N11264, N11290, N9775, N9769, N8902, N9899, N9975, N9626, N9685, N11296, N9149, N11183, N11231, N9971, N9565, N9560, N9276, N10886, N10888, N10331, N10330, N9896, N10329, N10328, N11002, N11004, N9103, N10028, AND3_3434_inw1, AND3_3436_inw1, AND3_3433_inw1, AND3_3435_inw1, N10439, N9561, N10026, N11106, N11108, N9557, N9758, N10264, N10002, N10961, N10963, N9220, N10205, N10204, N10203, N10773, N11073, N11075, N9344, N10598, N10344, N10265, N11267, N11269, N9385, N9375, N8966, N9715, N10771, N10659, N9206, N11298, N11297, N9223, N11185, N11187, N9995, N9596, N9591, N10895, N10897, N10866, N10340, N10339, N9892, N10338, N10337, N11011, N11013, N9165, N10766, N10024, AND3_3438_inw1, AND3_3440_inw1, AND3_3437_inw1, AND3_3439_inw1, N10444, N9592, N10765, N10023, N11110, N11112, N9791, N10719, N11342, N11302, OR4_3421_inw2, N11289, N11152, N11153, N10375, N10581, N10582, N10479, N10465, N11228, N11229, N10497, N10101, N10104, N8863, N7100, N9258, N9259, N7826, N8394, N9400, N9401, N9024, N9025, N7057, N8727, N8943, N9260, N9261, N8865, N8866, N8627, N8861, N9256, N9257, N10113, N9907, N10114, N9909, N8959, AND3_2232_inw1, g39_inw2, AND3_2080_inw1, N8992, AND3_2192_inw1, N8991, N9367, N9368, N10155, N9948, N9054, AND3_2252_inw1, N9053, N9417, N9418, N8811, N9615, AND3_2532_inw1, N9614, N8548, N9035, N9815, N9816, N8956, N8412, N9813, N9814, N9612, N9613, N8730, N8405, N10548, N9581, N9786, N8541, N9478, N9616, N9820, N9802, N9803, N9604, N9605, N9488, AND3_2530_inw1, N9603, AND3_2516_inw1, N9602, N9800, N9801, AND3_2518_inw1, N9485, N9624, AND3_2548_inw1, N9623, N9829, N9830, N9517, N9622, AND3_2546_inw1, N9621, N9827, N9828, N9520, N9690, N10953, N11006, N10531, N9835, N10838, N10103, n_352, N10021, n_317, N10014, N10649, N10648, n_332, N10017, N10296, N10391, N10367, N10354, N9543, N8857, N9072, N10729, N10170, N10317, N10316, N10566, N10431, N9071, N11299, N11288, N10432, N9077, N10180, N9093, N10057, AND3_2827_inw1, N10058, AND4_2861_inw2, g5_inw1, N10327, N10326, N10039, AND3_2834_inw1, N10040, AND4_2851_inw2, g75_inw1, N9551, N8871, N10557, N10437, N9092, N10438, N9098, N10762, N10321, N10248, N10555, N10318, N8881, N10761, N10708, N10760, N10707, OR4_2892_inw1, OR4_2906_inw1, N10535, N10534, N9935, N9575, N9897, N10750, N9978, N10621, N9695, N9768, N10528, N10440, N10525, N9563, N10042, N10060, AND3_2850_inw1, AND3_2860_inw1, AND4_2828_inw1, AND4_2835_inw1, N10341, N9721, N10652, N10545, N10544, N9949, N9608, N10769, N10626, N9720, N11317, N11309, N10627, N9726, N10907, N10539, N10445, N10767, N10536, N9594, N10906, N10865, N11227, N11226, N10905, N10864, OR3_2893_inw1, OR3_2907_inw1, N11312, N11315, N11205, OR4_3421_inw1, N10589, OR4_3183_inw2, OR4_3453_inw2, N9653, N8404, N10055, AND3_2830_inw1, N10056, AND4_2717_inw2, g34_inw1, N9698, N10050, N9323, OR4_2905_inw1, N9656, N10038, N9262, N9650, AND4_3022_inw1, AND4_3020_inw1, N9702, AND4_3023_inw1, N9727, N10067, N9412, N9408, N9618, N9617, N9986, N9585, N9582, N9332, N9983, N10231, N9324, N9326, N10704, N9733, N9402, N10232, N9784, N9785, AND3_2858_inw1, AND4_2831_inw1, N9992, N10238, N9806, N9989, N10237, N9805, N10007, N10239, N9825, N10010, N10240, N9826, N10690, N10689, OR4_3183_inw1, N10450, N10547, N10583, N10550, N9905, N10315, N10314, N10512, N10509, N11313, N11314, N10325, N10324, N10522, N9917, N10519, N10517, N10515, N10691, N10132, N10812, N10687, N10685, N10543, N10542, N10784, N10701, N10160, N10698, N11329, N11331, N10696, N10694, OR4_3453_inw1, N11327, N11320, N11246, N10739, N11257, N9908, N9939, N9938, N10134, N9911, N9910, N10115, N9906, N10399, N10388, N9947, N10402, N9954, N9953, N10161, N10138, N10137, N10136, N10135, N10293, N10629, N10294, N10159, N10158, N10300, N10157, N10156, N10299, N10163, N10162, N10306, N10165, N10164, N10307, N10673, N10671, N11328, N11321, N10683, N10681, N10815, N10890, N10825, N10823, N11338, N11335, N11333, N10836, N11286, AND3_3099_inw1, N10574, N10577, N10576, N10575, AND4_3020_inw2, AND4_3022_inw2, AND4_3023_inw2, N11334, N11340;
	assign N1490 = N1;
	assign N889 = N1;
	assign N388 = N1;
	assign N387 = N1;
	assign N1781 = ( N163 & N1 );
	assign N585 = ~N5;
	assign N628 = ~( N12 & N9 );
	assign N582 = ~N15;
	assign N1782 = ( N170 & N18 );
	assign N1793 = ( N169 & N18 );
	assign N1794 = ( N168 & N18 );
	assign N1795 = ( N167 & N18 );
	assign N1796 = ( N166 & N18 );
	assign N1797 = ( N165 & N18 );
	assign N1798 = ( N164 & N18 );
	assign N1811 = ( N177 & N18 );
	assign N1812 = ( N176 & N18 );
	assign N1813 = ( N175 & N18 );
	assign N1814 = ( N174 & N18 );
	assign N1815 = ( N173 & N18 );
	assign N1816 = ( N157 & N18 );
	assign N1817 = ( N156 & N18 );
	assign N1818 = ( N155 & N18 );
	assign N1819 = ( N154 & N18 );
	assign N1820 = ( N153 & N18 );
	assign N1857 = ( N181 & N18 );
	assign N1858 = ( N171 & N18 );
	assign N1859 = ( N180 & N18 );
	assign N1860 = ( N179 & N18 );
	assign N1861 = ( N178 & N18 );
	assign N1862 = ( N161 & N18 );
	assign N1863 = ( N151 & N18 );
	assign N1864 = ( N160 & N18 );
	assign N1865 = ( N159 & N18 );
	assign N1866 = ( N158 & N18 );
	assign N1957 = ( N209 & N18 );
	assign N1958 = ( N216 & N18 );
	assign N1959 = ( N215 & N18 );
	assign N1960 = ( N214 & N18 );
	assign N1961 = ( N213 & N18 );
	assign N1962 = ( N212 & N18 );
	assign N1963 = ( N211 & N18 );
	assign N1989 = ( N642 & N18 );
	assign N1990 = ( N644 & N18 );
	assign N1991 = ( N651 & N18 );
	assign N1992 = ( N674 & N18 );
	assign N1993 = ( N660 & N18 );
	assign N1994 = ( N666 & N18 );
	assign N1995 = ( N672 & N18 );
	assign N1996 = ( N673 & N18 );
	assign N2064 = ( N706 & N18 );
	assign N2065 = ( N708 & N18 );
	assign N2066 = ( N715 & N18 );
	assign N2067 = ( N721 & N18 );
	assign N2068 = ( N727 & N18 );
	assign N2069 = ( N599 & N18 );
	assign N2070 = ( N734 & N18 );
	assign N2071 = ( N742 & N18 );
	assign N2072 = ( N604 & N18 );
	assign N2073 = ( N609 & N18 );
	assign N2337 = ( N208 & N18 );
	assign N2338 = ( N198 & N18 );
	assign N2339 = ( N207 & N18 );
	assign N2340 = ( N206 & N18 );
	assign N2341 = ( N205 & N18 );
	assign N2374 = ( N193 & N18 );
	assign N2375 = ( N192 & N18 );
	assign N2376 = ( N191 & N18 );
	assign N2377 = ( N190 & N18 );
	assign N2378 = ( N189 & N18 );
	assign N2913 = ( N204 & N18 );
	assign N2914 = ( N203 & N18 );
	assign N2915 = ( N202 & N18 );
	assign N2916 = ( N201 & N18 );
	assign N2917 = ( N200 & N18 );
	assign N2918 = ( N235 & N18 );
	assign N2919 = ( N234 & N18 );
	assign N2920 = ( N233 & N18 );
	assign N2921 = ( N232 & N18 );
	assign N2922 = ( N231 & N18 );
	assign N2923 = ( N197 & N18 );
	assign N2924 = ( N187 & N18 );
	assign N2925 = ( N196 & N18 );
	assign N2926 = ( N195 & N18 );
	assign N2927 = ( N194 & N18 );
	assign N2928 = ( N227 & N18 );
	assign N2929 = ( N217 & N18 );
	assign N2930 = ( N226 & N18 );
	assign N2931 = ( N225 & N18 );
	assign N2932 = ( N224 & N18 );
	assign N2933 = ( N239 & N18 );
	assign N2934 = ( N229 & N18 );
	assign N2935 = ( N238 & N18 );
	assign N2936 = ( N237 & N18 );
	assign N2937 = ( N236 & N18 );
	assign N3005 = ( N223 & N18 );
	assign N3006 = ( N222 & N18 );
	assign N3007 = ( N221 & N18 );
	assign N3008 = ( N220 & N18 );
	assign N3009 = ( N219 & N18 );
	assign N3020 = ( N812 & N18 );
	assign N3021 = ( N814 & N18 );
	assign N3022 = ( N821 & N18 );
	assign N3023 = ( N827 & N18 );
	assign N3024 = ( N833 & N18 );
	assign N3025 = ( N839 & N18 );
	assign N3026 = ( N845 & N18 );
	assign N3027 = ( N853 & N18 );
	assign N3028 = ( N859 & N18 );
	assign N3029 = ( N865 & N18 );
	assign N3032 = ( N758 & N18 );
	assign N3033 = ( N759 & N18 );
	assign N3034 = ( N762 & N18 );
	assign N3035 = ( N768 & N18 );
	assign N3036 = ( N774 & N18 );
	assign N3037 = ( N780 & N18 );
	assign N3038 = ( N786 & N18 );
	assign N3039 = ( N794 & N18 );
	assign N3040 = ( N800 & N18 );
	assign N3041 = ( N806 & N18 );
	assign N695 = ~N18;
	assign N2674 = ( N2366 | N18 );
	assign N2680 = ( N2367 | N18 );
	assign N1930 = ( N23 & N695 );
	assign N1929 = ( N26 & N695 );
	assign N1928 = ( N29 & N695 );
	assign N2012 = ( N32 & N695 );
	assign N2011 = ( N35 & N695 );
	assign N1167 = ( N700 & N38 );
	assign N1537 = ( N957 & N38 );
	assign N1649 = ( N1029 & N38 );
	assign N1966 = ( N1222 & N38 );
	assign N2107 = ~( N38 & N1821 );
	assign N2268 = ~( N38 & N688 );
	assign N2355 = ~( N38 & N2171 );
	assign N2653 = ~( N38 & N1028 );
	assign N1708 = ~( N957 | N38 );
	assign N1822 = ~N38;
	assign N1927 = ( N41 & N695 );
	assign N1926 = ( N44 & N695 );
	assign N2010 = ( N47 & N695 );
	assign N2013 = ( N50 & N695 );
	assign N2424 = ( N53 & N695 );
	assign N2425 = ( N54 & N695 );
	assign N2426 = ( N55 & N695 );
	assign N2427 = ( N56 & N695 );
	assign N467 = ~N57;
	assign N2396 = ( N58 & N695 );
	assign N2399 = ( N59 & N695 );
	assign N2403 = ( N60 & N695 );
	assign N2404 = ( N61 & N695 );
	assign N2405 = ( N62 & N695 );
	assign N2434 = ( N63 & N695 );
	assign N2433 = ( N64 & N695 );
	assign N2429 = ( N65 & N695 );
	assign N2014 = ( N66 & N695 );
	assign N2418 = ( N69 & N695 );
	assign N2367 = ( N70 & N695 );
	assign N2423 = ( N73 & N695 );
	assign N2420 = ( N74 & N695 );
	assign N2422 = ( N75 & N695 );
	assign N2421 = ( N76 & N695 );
	assign N2397 = ( N77 & N695 );
	assign N2398 = ( N78 & N695 );
	assign N2402 = ( N79 & N695 );
	assign N2401 = ( N80 & N695 );
	assign N2400 = ( N81 & N695 );
	assign N2428 = ( N82 & N695 );
	assign N2430 = ( N83 & N695 );
	assign N2431 = ( N84 & N695 );
	assign N2432 = ( N85 & N695 );
	assign N2435 = ( N86 & N695 );
	assign N2361 = ( N87 & N695 );
	assign N2363 = ( N88 & N695 );
	assign AND4_2717_inw1 = ~( N89 & N9408 );
	assign N9407 = ~( N8548 & N89 );
	assign n_333 = ( N89 & N9408 );
	assign N2324 = ( N94 & N695 );
	assign N2323 = ( N97 & N695 );
	assign N2303 = ( N100 & N695 );
	assign N2299 = ( N103 & N695 );
	assign N945 = N106;
	assign N4467 = ~( N2632 & N106 );
	assign N674 = ~N106;
	assign N2436 = ( N109 & N695 );
	assign N2437 = ( N110 & N695 );
	assign N2360 = ( N111 & N695 );
	assign N2362 = ( N112 & N695 );
	assign N2359 = ( N113 & N695 );
	assign N2358 = ( N114 & N695 );
	assign N2321 = ( N115 & N695 );
	assign N2322 = ( N118 & N695 );
	assign N2325 = ( N121 & N695 );
	assign N2302 = ( N124 & N695 );
	assign N2301 = ( N127 & N695 );
	assign N2300 = ( N130 & N695 );
	assign N469 = ( N134 & N133 );
	assign N2281 = ( N135 & N695 );
	assign N2279 = ( N138 & N695 );
	assign N2277 = ( N141 & N695 );
	assign N2280 = ( N144 & N695 );
	assign N2278 = ( N147 & N695 );
	assign AND4_21_inw1 = ~( N150 & N184 );
	assign AND4_42_inw1 = ~( N210 & N152 );
	assign AND4_11_inw1 = ~( N162 & N172 );
	assign AND4_41_inw1 = ~( N183 & N182 );
	assign AND4_41_inw2 = ~( N185 & N186 );
	assign AND4_11_inw2 = ~( N188 & N199 );
	assign AND4_42_inw2 = ~( N218 & N230 );
	assign AND4_21_inw2 = ~( N228 & N240 );
	assign N1110 = ~( N242 & N585 );
	assign N2364 = ( N245 & N695 );
	assign N641 = ~N245;
	assign N478 = N248;
	assign N642 = ~N248;
	assign N643 = N251;
	assign N4471 = ~( N2619 & N251 );
	assign N644 = ~N251;
	assign N482 = N254;
	assign N4469 = ~( N2626 & N254 );
	assign N651 = ~N254;
	assign N484 = N257;
	assign N4465 = ~( N2638 & N257 );
	assign N660 = ~N257;
	assign N486 = N260;
	assign N4463 = ~( N2644 & N260 );
	assign N666 = ~N260;
	assign N489 = N263;
	assign N688 = ( N382 & N263 );
	assign N672 = ~N263;
	assign N492 = N267;
	assign N700 = ~( N382 & N267 );
	assign N673 = ~N267;
	assign N2365 = ( N271 & N695 );
	assign N705 = ~N271;
	assign N501 = N274;
	assign N706 = ~N274;
	assign N707 = N277;
	assign N4523 = ~( N2554 & N277 );
	assign N708 = ~N277;
	assign N505 = N280;
	assign N4519 = ~( N2561 & N280 );
	assign N715 = ~N280;
	assign N507 = N283;
	assign N4517 = ~( N2567 & N283 );
	assign N721 = ~N283;
	assign N509 = N286;
	assign N4515 = ~( N2573 & N286 );
	assign N727 = ~N286;
	assign N511 = N289;
	assign N4513 = ~( N2482 & N289 );
	assign N599 = ~N289;
	assign N513 = N293;
	assign N4521 = ~( N2488 & N293 );
	assign N734 = ~N293;
	assign N515 = N296;
	assign N4511 = ~( N2496 & N296 );
	assign N742 = ~N296;
	assign N517 = N299;
	assign N4509 = ~( N2502 & N299 );
	assign N604 = ~N299;
	assign N519 = N303;
	assign N4507 = ~( N2508 & N303 );
	assign N609 = ~N303;
	assign N535 = N307;
	assign N758 = ~N307;
	assign N537 = N310;
	assign N759 = ~N310;
	assign N539 = N313;
	assign N5958 = ~( N3343 & N313 );
	assign N762 = ~N313;
	assign N541 = N316;
	assign N5956 = ~( N3349 & N316 );
	assign N768 = ~N316;
	assign N543 = N319;
	assign N5954 = ~( N3355 & N319 );
	assign N774 = ~N319;
	assign N545 = N322;
	assign N5952 = ~( N3267 & N322 );
	assign N780 = ~N322;
	assign N547 = N325;
	assign N5950 = ~( N3273 & N325 );
	assign N786 = ~N325;
	assign N549 = N328;
	assign N5948 = ~( N3281 & N328 );
	assign N794 = ~N328;
	assign N551 = N331;
	assign N5946 = ~( N3287 & N331 );
	assign N800 = ~N331;
	assign N553 = N334;
	assign N5944 = ~( N3293 & N334 );
	assign N806 = ~N334;
	assign N556 = N337;
	assign N812 = ~N337;
	assign N813 = N340;
	assign N6076 = ~( N3315 & N340 );
	assign N814 = ~N340;
	assign N559 = N343;
	assign N6074 = ~( N3322 & N343 );
	assign N821 = ~N343;
	assign N561 = N346;
	assign N6072 = ~( N3328 & N346 );
	assign N827 = ~N346;
	assign N563 = N349;
	assign N6070 = ~( N3334 & N349 );
	assign N833 = ~N349;
	assign N565 = N352;
	assign N6068 = ~( N3384 & N352 );
	assign N839 = ~N352;
	assign N567 = N355;
	assign N6066 = ~( N3390 & N355 );
	assign N845 = ~N355;
	assign N569 = N358;
	assign N6064 = ~( N3398 & N358 );
	assign N853 = ~N358;
	assign N571 = N361;
	assign N6062 = ~( N3404 & N361 );
	assign N859 = ~N361;
	assign N573 = N364;
	assign N6060 = ~( N3410 & N364 );
	assign N865 = ~N364;
	assign N9288 = ( N367 & N8326 );
	assign N9767 = ( N9280 & N367 );
	assign N11316 = ( N367 & N11307 );
	assign AND3_2476_inw1 = ~( N367 & N8326 );
	assign AND3_2853_inw1 = ~( N367 & N9775 );
	assign AND3_2863_inw1 = ~( N367 & N9754 );
	assign N11224 = ~( AND3_3435_inw1 | N367 );
	assign N11225 = ~( AND3_3436_inw1 | N367 );
	assign AND4_2475_inw1 = ~( N367 & N8326 );
	assign AND4_2851_inw1 = ~( N367 & N9775 );
	assign AND4_2861_inw1 = ~( N367 & N9754 );
	assign N9773 = ~( N9307 & N367 );
	assign N9893 = ~( N367 & N9741 );
	assign N1115 = ~N367;
	assign n_318 = ( N367 & N9754 );
	assign n_353 = ( N367 & N9775 );
	assign N1028 = ( N382 & N641 );
	assign N1029 = ~( N382 & N705 );
	assign N241_O = N241_I;
	assign N1109 = ( N469 & N585 );
	assign N881 = ~( N467 & N585 );
	assign N2441 = ( N2239 & N628 );
	assign N2446 = ( N2241 & N628 );
	assign N2450 = ( N2242 & N628 );
	assign N2454 = ( N2243 & N628 );
	assign N2458 = ( N2244 & N628 );
	assign N2462 = ( N2247 & N628 );
	assign N2466 = ( N2248 & N628 );
	assign N2470 = ( N2249 & N628 );
	assign N2474 = ( N2250 & N628 );
	assign N2478 = ( N2251 & N628 );
	assign N2482 = ( N2252 & N628 );
	assign N2488 = ( N2253 & N628 );
	assign N2496 = ( N2254 & N628 );
	assign N2502 = ( N2255 & N628 );
	assign N2508 = ( N2256 & N628 );
	assign N2619 = ( N2348 & N628 );
	assign N2626 = ( N2349 & N628 );
	assign N2632 = ( N2350 & N628 );
	assign N2638 = ( N2351 & N628 );
	assign N2644 = ( N2352 & N628 );
	assign N2766 = ( N2354 & N628 );
	assign N2769 = ( N2353 & N628 );
	assign N2772 = ( N2246 & N628 );
	assign N2775 = ( N2245 & N628 );
	assign N4490 = ~( N2619 & N628 );
	assign N4496 = ~( N628 & N2441 );
	assign N5322 = ~( N628 & N4651 );
	assign N3073 = ~N628;
	assign g43_inw1 = ~( N628 & N6047 );
	assign N1114 = N582;
	assign N1111 = N582;
	assign N2239 = ( N695 | N1782 );
	assign N2241 = ( N695 | N1793 );
	assign N2242 = ( N695 | N1794 );
	assign N2243 = ( N695 | N1795 );
	assign N2244 = ( N695 | N1796 );
	assign N2245 = ( N695 | N1797 );
	assign N2246 = ( N695 | N1798 );
	assign N2247 = ( N695 | N1811 );
	assign N2248 = ( N695 | N1812 );
	assign N2249 = ( N695 | N1813 );
	assign N2250 = ( N695 | N1814 );
	assign N2251 = ( N695 | N1815 );
	assign N2252 = ( N695 | N1816 );
	assign N2253 = ( N695 | N1817 );
	assign N2254 = ( N695 | N1818 );
	assign N2255 = ( N695 | N1819 );
	assign N2256 = ( N695 | N1820 );
	assign N2793 = ( N2277 | N1857 );
	assign N2538 = ( N2278 | N1858 );
	assign N2542 = ( N2279 | N1859 );
	assign N2546 = ( N2280 | N1860 );
	assign N2550 = ( N2281 | N1861 );
	assign N2778 = ( N2277 | N1862 );
	assign N2554 = ( N2278 | N1863 );
	assign N2561 = ( N2279 | N1864 );
	assign N2567 = ( N2280 | N1865 );
	assign N2573 = ( N2281 | N1866 );
	assign N2348 = ( N695 | N1957 );
	assign N2349 = ( N695 | N1958 );
	assign N2350 = ( N695 | N1959 );
	assign N2351 = ( N695 | N1960 );
	assign N2352 = ( N695 | N1961 );
	assign N2353 = ( N695 | N1962 );
	assign N2354 = ( N695 | N1963 );
	assign N2781 = ( N2358 | N1989 );
	assign N2654 = ( N2359 | N1990 );
	assign N2658 = ( N2360 | N1991 );
	assign N2662 = ( N2361 | N1992 );
	assign N2666 = ( N2362 | N1993 );
	assign N2670 = ( N2363 | N1994 );
	assign N2787 = ( N2364 | N1995 );
	assign N2784 = ( N2365 | N1996 );
	assign N2796 = ( N2428 | N2064 );
	assign N2729 = ( N2429 | N2065 );
	assign N2733 = ( N2430 | N2066 );
	assign N2737 = ( N2431 | N2067 );
	assign N2741 = ( N2432 | N2068 );
	assign N2745 = ( N2433 | N2069 );
	assign N2749 = ( N2434 | N2070 );
	assign N2753 = ( N2435 | N2071 );
	assign N2757 = ( N2436 | N2072 );
	assign N2761 = ( N2437 | N2073 );
	assign N2790 = ( N2337 | N1926 );
	assign N2604 = ( N2338 | N1927 );
	assign N2607 = ( N2339 | N1928 );
	assign N2611 = ( N2340 | N1929 );
	assign N2615 = ( N2341 | N1930 );
	assign N2688 = ( N2374 | N2010 );
	assign N2692 = ( N2375 | N2011 );
	assign N2696 = ( N2376 | N2012 );
	assign N2700 = ( N2377 | N2013 );
	assign N2704 = ( N2378 | N2014 );
	assign N3247 = ( N2913 | N2299 );
	assign N3251 = ( N2914 | N2300 );
	assign N3255 = ( N2915 | N2301 );
	assign N3259 = ( N2916 | N2302 );
	assign N3263 = ( N2917 | N2303 );
	assign N3267 = ( N2918 | N2299 );
	assign N3273 = ( N2919 | N2300 );
	assign N3281 = ( N2920 | N2301 );
	assign N3287 = ( N2921 | N2302 );
	assign N3293 = ( N2922 | N2303 );
	assign N3789 = ( N2923 | N2321 );
	assign N3299 = ( N2924 | N2322 );
	assign N3303 = ( N2925 | N2323 );
	assign N3307 = ( N2926 | N2324 );
	assign N3311 = ( N2927 | N2325 );
	assign N3783 = ( N2928 | N2321 );
	assign N3315 = ( N2929 | N2322 );
	assign N3322 = ( N2930 | N2323 );
	assign N3328 = ( N2931 | N2324 );
	assign N3334 = ( N2932 | N2325 );
	assign N3786 = ( N2933 | N1926 );
	assign N3340 = ( N2934 | N1927 );
	assign N3343 = ( N2935 | N1928 );
	assign N3349 = ( N2936 | N1929 );
	assign N3355 = ( N2937 | N1930 );
	assign N3384 = ( N3005 | N2010 );
	assign N3390 = ( N3006 | N2011 );
	assign N3398 = ( N3007 | N2012 );
	assign N3404 = ( N3008 | N2013 );
	assign N3410 = ( N3009 | N2014 );
	assign N3891 = ( N3020 | N2396 );
	assign N3416 = ( N3021 | N2397 );
	assign N3420 = ( N3022 | N2398 );
	assign N3424 = ( N3023 | N2399 );
	assign N3428 = ( N3024 | N2400 );
	assign N3432 = ( N3025 | N2401 );
	assign N3436 = ( N3026 | N2402 );
	assign N3440 = ( N3027 | N2403 );
	assign N3444 = ( N3028 | N2404 );
	assign N3448 = ( N3029 | N2405 );
	assign N3888 = ( N3032 | N2418 );
	assign N3885 = ( N3033 | N2367 );
	assign N3454 = ( N3034 | N2420 );
	assign N3458 = ( N3035 | N2421 );
	assign N3462 = ( N3036 | N2422 );
	assign N3466 = ( N3037 | N2423 );
	assign N3470 = ( N3038 | N2424 );
	assign N3474 = ( N3039 | N2425 );
	assign N3478 = ( N3040 | N2426 );
	assign N3482 = ( N3041 | N2427 );
	assign N2366 = ( N759 & N695 );
	assign N3381 = ( N695 & N2604 );
	assign N4769 = ( N3340 & N695 );
	assign N5960 = ( N2674 & N4769 );
	assign N7744 = ~( N2674 & N6968 );
	assign N6217 = ~( N2674 | N4769 );
	assign N4575 = ~N2674;
	assign N6690 = ~( N2680 & N6165 );
	assign N4768 = ~N2680;
	assign n_350 = ( N7358 & N2680 );
	assign N3507 = ~( N1167 | N2866 );
	assign OR3_922_inw1 = ~( N1167 | N2866 );
	assign N2866 = ( N2257 & N1537 );
	assign N4488 = ~( N1537 & N3954 );
	assign N6712 = ~( N1537 & N3126 );
	assign N2537 = ~N1537;
	assign N4193 = ( N1649 | N3379 );
	assign N3379 = ( N2650 & N1966 );
	assign N2257 = ~( N2107 & N2108 );
	assign N2523 = ~( N2268 & N2111 );
	assign N2650 = ~( N2355 & N2172 );
	assign N2988 = ~( N2653 & N2357 );
	assign N4487 = ~( N1708 & N3954 );
	assign N6711 = ~( N1708 & N6191 );
	assign N2117 = ~N1708;
	assign N2108 = ~( N700 & N1822 );
	assign N2111 = ~( N957 & N1822 );
	assign N2172 = ~( N1029 & N1822 );
	assign N2357 = ~( N1222 & N1822 );
	assign N9790 = ~( AND4_2717_inw1 | AND4_2717_inw2 );
	assign N9817 = ( N9617 & N9407 );
	assign g34_inw2 = ~( N8421 & n_333 );
	assign N5654 = ~( N4467 & N5169 );
	assign N3101 = ( N674 & N2632 );
	assign N5169 = ~( N674 & N4468 );
	assign N528 = ~( AND4_21_inw1 | AND4_21_inw2 );
	assign N578 = ~( AND4_42_inw1 | AND4_42_inw2 );
	assign N494 = ~( AND4_11_inw1 | AND4_11_inw2 );
	assign N575 = ~( AND4_41_inw1 | AND4_41_inw2 );
	assign N1112 = N1110;
	assign N5683 = ~( N4471 & N5171 );
	assign N3114 = ( N644 & N2619 );
	assign N5171 = ~( N644 & N4472 );
	assign N3515 = ~( N644 | N2619 );
	assign N5670 = ~( N4469 & N5170 );
	assign N3107 = ( N651 & N2626 );
	assign N5170 = ~( N651 & N4470 );
	assign N5640 = ~( N4465 & N5168 );
	assign N3097 = ( N660 & N2638 );
	assign N5168 = ~( N660 & N4466 );
	assign N5632 = ~( N4463 & N5167 );
	assign N3096 = ( N666 & N2644 );
	assign N5167 = ~( N666 & N4464 );
	assign N957 = ~N688;
	assign N1821 = ~N700;
	assign N5856 = ~( N4523 & N5204 );
	assign N3202 = ( N708 & N2554 );
	assign N5204 = ~( N708 & N4501 );
	assign N3628 = ~( N708 | N2554 );
	assign N5837 = ~( N4519 & N5202 );
	assign N3195 = ( N715 & N2561 );
	assign N5202 = ~( N715 & N4504 );
	assign N5821 = ~( N4517 & N5201 );
	assign N3189 = ( N721 & N2567 );
	assign N5201 = ~( N721 & N4503 );
	assign N5807 = ~( N4515 & N5200 );
	assign N3185 = ( N727 & N2573 );
	assign N5200 = ~( N727 & N4506 );
	assign N5799 = ~( N4513 & N5199 );
	assign N3184 = ( N599 & N2482 );
	assign N5199 = ~( N599 & N4505 );
	assign N5850 = ~( N4521 & N5203 );
	assign N3178 = ( N734 & N2488 );
	assign N5203 = ~( N734 & N4522 );
	assign N3625 = ~( N734 | N2488 );
	assign N5789 = ~( N4511 & N5198 );
	assign N3173 = ( N742 & N2496 );
	assign N5198 = ~( N742 & N4512 );
	assign N5778 = ~( N4509 & N5197 );
	assign N3169 = ( N604 & N2502 );
	assign N5197 = ~( N604 & N4510 );
	assign N5771 = ~( N4507 & N5196 );
	assign N3168 = ( N609 & N2508 );
	assign N5196 = ~( N609 & N4508 );
	assign N6957 = ~( N5958 & N6547 );
	assign N4570 = ( N762 & N3343 );
	assign N6547 = ~( N762 & N5959 );
	assign N6946 = ~( N5956 & N6546 );
	assign N4566 = ( N768 & N3349 );
	assign N6546 = ~( N768 & N5957 );
	assign N6936 = ~( N5954 & N6545 );
	assign N4563 = ( N774 & N3355 );
	assign N6545 = ~( N774 & N5955 );
	assign N6929 = ~( N5952 & N6544 );
	assign N4562 = ( N780 & N3267 );
	assign N6544 = ~( N780 & N5953 );
	assign N6923 = ~( N5950 & N6543 );
	assign N4555 = ( N3273 & N786 );
	assign N6543 = ~( N786 & N5951 );
	assign N4844 = ~( N3273 | N786 );
	assign N6912 = ~( N5948 & N6542 );
	assign N4549 = ( N794 & N3281 );
	assign N6542 = ~( N794 & N5949 );
	assign N6901 = ~( N5946 & N6541 );
	assign N4545 = ( N800 & N3287 );
	assign N6541 = ~( N800 & N5947 );
	assign N6894 = ~( N5944 & N6540 );
	assign N4544 = ( N806 & N3293 );
	assign N6540 = ~( N806 & N5945 );
	assign N7180 = ~( N6076 & N6629 );
	assign N4687 = ( N814 & N3315 );
	assign N6629 = ~( N814 & N6077 );
	assign N5030 = ~( N814 | N3315 );
	assign N7170 = ~( N6074 & N6628 );
	assign N4682 = ( N821 & N3322 );
	assign N6628 = ~( N821 & N6075 );
	assign N7159 = ~( N6072 & N6627 );
	assign N4678 = ( N827 & N3328 );
	assign N6627 = ~( N827 & N6073 );
	assign N7149 = ~( N6070 & N6626 );
	assign N4675 = ( N833 & N3334 );
	assign N6626 = ~( N833 & N6071 );
	assign N7142 = ~( N6068 & N6625 );
	assign N4674 = ( N839 & N3384 );
	assign N6625 = ~( N839 & N6069 );
	assign N7136 = ~( N6066 & N6624 );
	assign N4667 = ( N3390 & N845 );
	assign N6624 = ~( N845 & N6067 );
	assign N4940 = ~( N3390 | N845 );
	assign N7125 = ~( N6064 & N6623 );
	assign N4661 = ( N853 & N3398 );
	assign N6623 = ~( N853 & N6065 );
	assign N7114 = ~( N6062 & N6622 );
	assign N4657 = ( N859 & N3404 );
	assign N6622 = ~( N859 & N6063 );
	assign N7107 = ~( N6060 & N6621 );
	assign N4656 = ( N865 & N3410 );
	assign N6621 = ~( N865 & N6061 );
	assign N9635 = ( N5960 | N9288 );
	assign g87_inw2 = ~( N6936 & N9288 );
	assign N9925 = ( N8902 | N9767 );
	assign N11323 = ( N11308 | N11316 );
	assign N9287 = ~( AND3_2476_inw1 | N6957 );
	assign N10043 = ~( AND3_2853_inw1 | N9385 );
	assign N10061 = ~( AND3_2863_inw1 | N9344 );
	assign OR4_3452_inw2 = ~( N11224 | N11225 );
	assign N9286 = ~( AND4_2475_inw1 | AND4_2475_inw2 );
	assign N10041 = ~( AND4_2851_inw1 | AND4_2851_inw2 );
	assign N10059 = ~( AND4_2861_inw1 | AND4_2861_inw2 );
	assign N9932 = ( N9575 & N9773 );
	assign N10025 = ~( N9740 & N9893 );
	assign N11308 = ( N11296 & N1115 );
	assign N11222 = ~( AND3_3433_inw1 | N1115 );
	assign N11223 = ~( AND3_3434_inw1 | N1115 );
	assign N9740 = ~( N8326 & N1115 );
	assign g5_inw2 = ~( N8269 & n_318 );
	assign g75_inw2 = ~( N8262 & n_353 );
	assign N1222 = ~N1028;
	assign N2171 = ~N1029;
	assign N1113 = ~N1109;
	assign N3080 = ~N2441;
	assign N3373 = ( N2658 & N2446 );
	assign N5185 = ~( N2446 & N4497 );
	assign N5320 = ~( N2446 & N4649 );
	assign N4498 = ~N2446;
	assign N5186 = ~( N2450 & N4498 );
	assign N5318 = ~( N2450 & N4647 );
	assign N4497 = ~N2450;
	assign g40_inw2 = ~( N2662 & N2450 );
	assign N3371 = ( N2666 & N2454 );
	assign N5187 = ~( N2454 & N4499 );
	assign N5316 = ~( N2454 & N4645 );
	assign N4500 = ~N2454;
	assign N3370 = ( N2670 & N2458 );
	assign N5188 = ~( N2458 & N4500 );
	assign N5314 = ~( N2458 & N4643 );
	assign N4499 = ~N2458;
	assign N3365 = ( N2745 & N2462 );
	assign N5289 = ~( N2462 & N4617 );
	assign N5433 = ~( N2462 & N4620 );
	assign N4618 = ~N2462;
	assign N3364 = ( N2749 & N2466 );
	assign N5297 = ~( N2466 & N4625 );
	assign N5584 = ~( N2466 & N4616 );
	assign N4626 = ~N2466;
	assign N5287 = ~( N2470 & N4615 );
	assign N5585 = ~( N2470 & N4626 );
	assign N4616 = ~N2470;
	assign g44_inw2 = ~( N2753 & N2470 );
	assign N3362 = ( N2757 & N2474 );
	assign N5285 = ~( N2474 & N4613 );
	assign N5586 = ~( N2474 & N4612 );
	assign N4614 = ~N2474;
	assign N3361 = ( N2761 & N2478 );
	assign N5283 = ~( N2478 & N4611 );
	assign N5587 = ~( N2478 & N4614 );
	assign N4612 = ~N2478;
	assign N5193 = ~( N2482 & N4506 );
	assign N4505 = ~N2482;
	assign N5474 = ~( N2488 & N4512 );
	assign N4522 = ~N2488;
	assign N5475 = ~( N2496 & N4522 );
	assign N4512 = ~N2496;
	assign N5476 = ~( N2502 & N4508 );
	assign N4510 = ~N2502;
	assign N5477 = ~( N2508 & N4510 );
	assign N4508 = ~N2508;
	assign N4472 = ~N2619;
	assign N5180 = ~( N2626 & N4468 );
	assign N4470 = ~N2626;
	assign N5181 = ~( N2632 & N4470 );
	assign N4468 = ~N2632;
	assign N5182 = ~( N2638 & N4464 );
	assign N4466 = ~N2638;
	assign N5183 = ~( N2644 & N4466 );
	assign N4464 = ~N2644;
	assign N4327 = ~( N2766 & N3552 );
	assign N3551 = ~N2766;
	assign N4326 = ~( N2769 & N3551 );
	assign N3552 = ~N2769;
	assign N4334 = ~( N2772 & N3570 );
	assign N3569 = ~N2772;
	assign N4333 = ~( N2775 & N3569 );
	assign N3570 = ~N2775;
	assign N5736 = ~( N5179 & N4490 );
	assign N5747 = ~( N5184 & N4496 );
	assign N6059 = ~( N5322 & N5323 );
	assign N5179 = ~( N3073 & N4472 );
	assign N5184 = ~( N3080 & N3073 );
	assign N5323 = ~( N2654 & N3073 );
	assign N7106 = ~( g43_inw1 | g43_inw2 );
	assign N5429 = ~( N2793 & N4628 );
	assign N3453 = ~N2793;
	assign N4751 = ~( N2538 & N3453 );
	assign N5299 = ~( N2538 & N4627 );
	assign N4628 = ~N2538;
	assign g62_inw1 = ~( N2538 & N6009 );
	assign N3368 = ( N2733 & N2542 );
	assign N5295 = ~( N2542 & N4623 );
	assign N5430 = ~( N2542 & N4622 );
	assign N4624 = ~N2542;
	assign N5293 = ~( N2546 & N4621 );
	assign N5431 = ~( N2546 & N4624 );
	assign N4622 = ~N2546;
	assign g59_inw2 = ~( N2737 & N2546 );
	assign N3366 = ( N2741 & N2550 );
	assign N5291 = ~( N2550 & N4619 );
	assign N5432 = ~( N2550 & N4618 );
	assign N4620 = ~N2550;
	assign N5189 = ~( N2778 & N4501 );
	assign N3167 = ~N2778;
	assign N4502 = ~( N2554 & N3167 );
	assign N4501 = ~N2554;
	assign N5190 = ~( N2561 & N4503 );
	assign N4504 = ~N2561;
	assign N5191 = ~( N2567 & N4504 );
	assign N4503 = ~N2567;
	assign N5192 = ~( N2573 & N4505 );
	assign N4506 = ~N2573;
	assign N5363 = ~( N2781 & N4651 );
	assign N3380 = ~N2781;
	assign N4694 = ~( N2654 & N3380 );
	assign N4651 = ~N2654;
	assign n_338 = ( N6041 & N2654 );
	assign N5321 = ~( N2658 & N4498 );
	assign N5364 = ~( N2658 & N4647 );
	assign N4649 = ~N2658;
	assign N5319 = ~( N2662 & N4497 );
	assign N5365 = ~( N2662 & N4649 );
	assign N4647 = ~N2662;
	assign N5317 = ~( N2666 & N4500 );
	assign N5366 = ~( N2666 & N4643 );
	assign N4645 = ~N2666;
	assign N5315 = ~( N2670 & N4499 );
	assign N5367 = ~( N2670 & N4645 );
	assign N4643 = ~N2670;
	assign N4411 = ~( N2787 & N3781 );
	assign N3782 = ~N2787;
	assign N4412 = ~( N2784 & N3782 );
	assign N3781 = ~N2784;
	assign N5451 = ~( N2796 & N4627 );
	assign N3486 = ~N2796;
	assign N4776 = ~( N2729 & N3486 );
	assign N5300 = ~( N2729 & N4628 );
	assign N4627 = ~N2729;
	assign n_346 = ( N6003 & N2729 );
	assign N5296 = ~( N2733 & N4624 );
	assign N5452 = ~( N2733 & N4621 );
	assign N4623 = ~N2733;
	assign N5294 = ~( N2737 & N4622 );
	assign N5453 = ~( N2737 & N4623 );
	assign N4621 = ~N2737;
	assign N5292 = ~( N2741 & N4620 );
	assign N5454 = ~( N2741 & N4617 );
	assign N4619 = ~N2741;
	assign N5290 = ~( N2745 & N4618 );
	assign N5455 = ~( N2745 & N4619 );
	assign N4617 = ~N2745;
	assign N5298 = ~( N2749 & N4626 );
	assign N5602 = ~( N2749 & N4615 );
	assign N4625 = ~N2749;
	assign N5288 = ~( N2753 & N4616 );
	assign N5603 = ~( N2753 & N4625 );
	assign N4615 = ~N2753;
	assign N5286 = ~( N2757 & N4614 );
	assign N5604 = ~( N2757 & N4611 );
	assign N4613 = ~N2757;
	assign N5284 = ~( N2761 & N4612 );
	assign N5605 = ~( N2761 & N4613 );
	assign N4611 = ~N2761;
	assign N5425 = ~( N2790 & N4745 );
	assign N3452 = ~N2790;
	assign N4746 = ~( N2604 & N3452 );
	assign N4745 = ~N2604;
	assign N4766 = ( N3454 & N2607 );
	assign N5426 = ~( N2607 & N4747 );
	assign N6687 = ~( N2607 & N6160 );
	assign N4748 = ~N2607;
	assign N5427 = ~( N2611 & N4748 );
	assign N6686 = ~( N2611 & N6158 );
	assign N4747 = ~N2611;
	assign g67_inw2 = ~( N3458 & N2611 );
	assign N4762 = ( N3462 & N2615 );
	assign N6668 = ~( N2615 & N6135 );
	assign N6685 = ~( N2615 & N6156 );
	assign N4749 = ~N2615;
	assign N4637 = ( N3432 & N2688 );
	assign N6597 = ~( N2688 & N6029 );
	assign N6661 = ~( N2688 & N6032 );
	assign N4636 = ~N2688;
	assign N4635 = ( N3436 & N2692 );
	assign N5571 = ~( N2692 & N4633 );
	assign N6604 = ~( N2692 & N6037 );
	assign N4642 = ~N2692;
	assign N5572 = ~( N2696 & N4642 );
	assign N6596 = ~( N2696 & N6027 );
	assign N4633 = ~N2696;
	assign g53_inw2 = ~( N3440 & N2696 );
	assign N4632 = ( N3444 & N2700 );
	assign N5573 = ~( N2700 & N4629 );
	assign N6595 = ~( N2700 & N6025 );
	assign N4631 = ~N2700;
	assign N4630 = ( N3448 & N2704 );
	assign N5574 = ~( N2704 & N4631 );
	assign N6594 = ~( N2704 & N6023 );
	assign N4629 = ~N2704;
	assign N4760 = ( N3466 & N3247 );
	assign N6136 = ~( N3247 & N4749 );
	assign N6683 = ~( N3247 & N6154 );
	assign N6135 = ~N3247;
	assign N4759 = ( N3470 & N3251 );
	assign N6688 = ~( N3251 & N6162 );
	assign N6741 = ~( N3251 & N6153 );
	assign N6163 = ~N3251;
	assign N6681 = ~( N3255 & N6152 );
	assign N6742 = ~( N3255 & N6163 );
	assign N6153 = ~N3255;
	assign g56_inw2 = ~( N3474 & N3255 );
	assign N4757 = ( N3478 & N3259 );
	assign N6679 = ~( N3259 & N6150 );
	assign N6743 = ~( N3259 & N6149 );
	assign N6151 = ~N3259;
	assign N4756 = ( N3482 & N3263 );
	assign N6677 = ~( N3263 & N6148 );
	assign N6744 = ~( N3263 & N6151 );
	assign N6149 = ~N3263;
	assign N6648 = ~( N3267 & N5955 );
	assign N5953 = ~N3267;
	assign N6733 = ~( N3273 & N5949 );
	assign N5951 = ~N3273;
	assign N6734 = ~( N3281 & N5951 );
	assign N5949 = ~N3281;
	assign N6735 = ~( N3287 & N5945 );
	assign N5947 = ~N3287;
	assign N6736 = ~( N3293 & N5947 );
	assign N5945 = ~N3293;
	assign N6658 = ~( N3789 & N6040 );
	assign N4743 = ~N3789;
	assign N6122 = ~( N3299 & N4743 );
	assign N6605 = ~( N3299 & N6039 );
	assign N6040 = ~N3299;
	assign g66_inw1 = ~( N3299 & N7086 );
	assign N4640 = ( N3420 & N3303 );
	assign N6602 = ~( N3303 & N6035 );
	assign N6659 = ~( N3303 & N6034 );
	assign N6036 = ~N3303;
	assign N6600 = ~( N3307 & N6033 );
	assign N6660 = ~( N3307 & N6036 );
	assign N6034 = ~N3307;
	assign g63_inw2 = ~( N3424 & N3307 );
	assign N4638 = ( N3428 & N3311 );
	assign N6125 = ~( N3311 & N4636 );
	assign N6598 = ~( N3311 & N6031 );
	assign N6032 = ~N3311;
	assign N6639 = ~( N3783 & N6077 );
	assign N4699 = ~N3783;
	assign N6091 = ~( N3315 & N4699 );
	assign N6077 = ~N3315;
	assign N6640 = ~( N3322 & N6073 );
	assign N6075 = ~N3322;
	assign N6641 = ~( N3328 & N6075 );
	assign N6073 = ~N3328;
	assign N6642 = ~( N3334 & N6069 );
	assign N6071 = ~N3334;
	assign N6644 = ~( N3786 & N6096 );
	assign N4700 = ~N3786;
	assign N6097 = ~( N3340 & N4700 );
	assign N6096 = ~N3340;
	assign N6645 = ~( N3343 & N5957 );
	assign N5959 = ~N3343;
	assign N6646 = ~( N3349 & N5959 );
	assign N5957 = ~N3349;
	assign N6647 = ~( N3355 & N5953 );
	assign N5955 = ~N3355;
	assign N6643 = ~( N3384 & N6071 );
	assign N6069 = ~N3384;
	assign N6729 = ~( N3390 & N6065 );
	assign N6067 = ~N3390;
	assign N6730 = ~( N3398 & N6067 );
	assign N6065 = ~N3398;
	assign N6731 = ~( N3404 & N6061 );
	assign N6063 = ~N3404;
	assign N6732 = ~( N3410 & N6063 );
	assign N6061 = ~N3410;
	assign N6706 = ~( N3891 & N6039 );
	assign N4783 = ~N3891;
	assign N6186 = ~( N3416 & N4783 );
	assign N6606 = ~( N3416 & N6040 );
	assign N6039 = ~N3416;
	assign n_348 = ( N7080 & N3416 );
	assign N6603 = ~( N3420 & N6036 );
	assign N6707 = ~( N3420 & N6033 );
	assign N6035 = ~N3420;
	assign N6601 = ~( N3424 & N6034 );
	assign N6708 = ~( N3424 & N6035 );
	assign N6033 = ~N3424;
	assign N6599 = ~( N3428 & N6032 );
	assign N6709 = ~( N3428 & N6029 );
	assign N6031 = ~N3428;
	assign N6030 = ~( N3432 & N4636 );
	assign N6710 = ~( N3432 & N6031 );
	assign N6029 = ~N3432;
	assign N6038 = ~( N3436 & N4642 );
	assign N6755 = ~( N3436 & N6027 );
	assign N6037 = ~N3436;
	assign N6028 = ~( N3440 & N4633 );
	assign N6756 = ~( N3440 & N6037 );
	assign N6027 = ~N3440;
	assign N6026 = ~( N3444 & N4631 );
	assign N6757 = ~( N3444 & N6023 );
	assign N6025 = ~N3444;
	assign N6024 = ~( N3448 & N4629 );
	assign N6758 = ~( N3448 & N6025 );
	assign N6023 = ~N3448;
	assign N5456 = ~( N3888 & N4781 );
	assign N4782 = ~N3888;
	assign N5457 = ~( N3885 & N4782 );
	assign N4781 = ~N3885;
	assign N6161 = ~( N3454 & N4748 );
	assign N6702 = ~( N3454 & N6158 );
	assign N6160 = ~N3454;
	assign N6159 = ~( N3458 & N4747 );
	assign N6703 = ~( N3458 & N6160 );
	assign N6158 = ~N3458;
	assign N6157 = ~( N3462 & N4749 );
	assign N6704 = ~( N3462 & N6154 );
	assign N6156 = ~N3462;
	assign N6684 = ~( N3466 & N6135 );
	assign N6705 = ~( N3466 & N6156 );
	assign N6154 = ~N3466;
	assign N6689 = ~( N3470 & N6163 );
	assign N6751 = ~( N3470 & N6152 );
	assign N6162 = ~N3470;
	assign N6682 = ~( N3474 & N6153 );
	assign N6752 = ~( N3474 & N6162 );
	assign N6152 = ~N3474;
	assign N6680 = ~( N3478 & N6151 );
	assign N6753 = ~( N3478 & N6148 );
	assign N6150 = ~N3478;
	assign N6678 = ~( N3482 & N6149 );
	assign N6754 = ~( N3482 & N6150 );
	assign N6148 = ~N3482;
	assign N6164 = ~( N3381 & N4768 );
	assign N6165 = ~N3381;
	assign g70_inw1 = ~( N3381 & N7364 );
	assign N6967 = ~( N4769 & N4575 );
	assign N6968 = ~N4769;
	assign N8357 = ( N6957 & N5960 );
	assign N8356 = ~( AND3_2117_inw1 | N5960 );
	assign AND4_2115_inw2 = ~( N5960 & N6936 );
	assign N9863 = ~( N5960 & N9690 );
	assign N8717 = ~N5960;
	assign g29_inw1 = ~( N6929 & N5960 );
	assign N8326 = ~( N6967 & N7744 );
	assign N10086 = ~( N6217 & N9975 );
	assign N7552 = ~N6217;
	assign N7377 = ~( N6164 & N6690 );
	assign g70_inw2 = ~( n_349 & n_350 );
	assign N5165 = ~( N3507 & N4473 );
	assign N6194 = ~( N3507 & N2537 );
	assign N9065 = ~( N3507 & N8609 );
	assign N3126 = ~N3507;
	assign N4303 = ~( OR3_922_inw1 & N3122 );
	assign N5178 = ~( N3955 & N4488 );
	assign N7444 = ~( N6194 & N6712 );
	assign N3955 = ~( N2257 & N2537 );
	assign N10451 = ( N10296 & N4193 );
	assign N5324 = ~N4193;
	assign n_331 = ( N4193 | N8960 );
	assign N3122 = ( N2523 & N2257 );
	assign N3953 = ~( N2257 & N2117 );
	assign N10271 = ~( N2257 & N10241 );
	assign N10272 = ~( N2257 & N10242 );
	assign N3954 = ~N2257;
	assign N10731 = ( N2523 & N10583 );
	assign N9955 = ~( N2523 & N9835 );
	assign N9956 = ~( N2523 & N9837 );
	assign N3135 = ~N2523;
	assign N3375 = ( N2988 & N2650 );
	assign N5177 = ~( N3953 & N4487 );
	assign N7441 = ~( N6192 & N6711 );
	assign N6192 = ~( N4784 & N2117 );
	assign OR4_2905_inw2 = ~( N10056 | N9790 );
	assign N10054 = ( N9817 & N9029 );
	assign N10053 = ~N9817;
	assign N9734 = ~( g34_inw1 | g34_inw2 );
	assign N6777 = ( N5654 & N3107 );
	assign AND3_1756_inw1 = ~( N5654 & N3107 );
	assign AND3_1763_inw1 = ~( N5670 & N5654 );
	assign AND3_1764_inw1 = ~( N5683 & N5654 );
	assign AND4_1753_inw1 = ~( N5654 & N5632 );
	assign AND4_1757_inw1 = ~( N5670 & N5654 );
	assign AND4_1758_inw1 = ~( N5683 & N5654 );
	assign AND4_2965_inw2 = ~( N5654 & N5670 );
	assign N10644 = ~( N5654 & N10570 );
	assign N11141 = ~( N5654 & N11114 );
	assign N11142 = ~( N5654 & N11116 );
	assign N8250 = ~N5654;
	assign n_320 = ( N5670 & N5654 );
	assign g11_inw1 = ~( N5654 & N5632 );
	assign g77_inw1 = ~( N5654 & N5640 );
	assign g95_inw1 = ~( N5654 & N5670 );
	assign N6770 = ( N5640 & N3101 );
	assign N6767 = ~( AND3_1752_inw1 | N3101 );
	assign NOR3_2032_inw1 = ~( N3101 | N6777 );
	assign OR4_2030_inw1 = ~( N3101 | N6777 );
	assign OR4_3029_inw1 = ~( N3101 | N6777 );
	assign N886 = ( N528 & N578 );
	assign N882 = ~N528;
	assign N883 = ~N578;
	assign N887 = ( N575 & N494 );
	assign N885 = ~N494;
	assign N884 = ~N575;
	assign N6783 = ( N5683 & N5670 );
	assign N10281 = ( N10141 & N5683 );
	assign AND3_2966_inw1 = ~( N10141 & N5683 );
	assign AND4_2965_inw1 = ~( N10141 & N5683 );
	assign N10565 = ~( N5683 & N10465 );
	assign N10737 = ~( N5683 & N10671 );
	assign N10738 = ~( N5683 & N10673 );
	assign N8247 = ~N5683;
	assign n_321 = ( N5640 & N5683 );
	assign N6782 = ( N5670 & N3114 );
	assign N6778 = ~( AND3_1763_inw1 | N3114 );
	assign AND4_1757_inw2 = ~( N3114 & N5640 );
	assign N9435 = ~( N3114 & N9072 );
	assign N6195 = ~N3114;
	assign N10428 = ( N3114 | N10281 );
	assign g9_inw1 = ~( N5632 & N3114 );
	assign N9432 = ~( N3515 & N9066 );
	assign N4795 = ~N3515;
	assign N6779 = ~( AND3_1764_inw1 | N5670 );
	assign N10280 = ~( AND3_2966_inw1 | N5670 );
	assign AND4_1758_inw2 = ~( N5640 & N5670 );
	assign N10645 = ~( N5670 & N10572 );
	assign N10909 = ~( N5670 & N10872 );
	assign N10910 = ~( N5670 & N10874 );
	assign N8251 = ~N5670;
	assign g11_inw2 = ~( N5670 & n_321 );
	assign AND4_1753_inw2 = ~( N3107 & N5640 );
	assign N7613 = ( N3107 | N6782 );
	assign OR3_3030_inw1 = ~( N3107 | N6782 );
	assign AND3_1752_inw1 = ~( N5640 & N5632 );
	assign N6771 = ~( AND3_1756_inw1 | N5640 );
	assign N10643 = ~( N5640 & N10568 );
	assign N11242 = ~( N5640 & N11213 );
	assign N11243 = ~( N5640 & N11215 );
	assign N8249 = ~N5640;
	assign g9_inw2 = ~( N5640 & n_320 );
	assign g95_inw2 = ~( N5640 & N10281 );
	assign N6766 = ( N5632 & N3097 );
	assign NOR4_2033_inw1 = ~( N3097 | N6770 );
	assign n_362 = ( N3097 | N6770 );
	assign N10642 = ~( N5632 & N10566 );
	assign N11023 = ~( N5632 & N10988 );
	assign N11024 = ~( N5632 & N10990 );
	assign N8248 = ~N5632;
	assign g77_inw2 = ~( N5632 & N6783 );
	assign n_319 = ( N3096 | N6766 );
	assign N6866 = ( N5856 & N5837 );
	assign N10290 = ( N10148 & N5856 );
	assign AND3_1816_inw1 = ~( N5856 & N5821 );
	assign AND3_2972_inw1 = ~( N10148 & N5856 );
	assign AND4_1810_inw1 = ~( N5856 & N5821 );
	assign AND4_2971_inw1 = ~( N10148 & N5856 );
	assign N10552 = ~( N5856 & N10455 );
	assign N10746 = ~( N5856 & N10681 );
	assign N10747 = ~( N5856 & N10683 );
	assign N8242 = ~N5856;
	assign n_322 = ( N5807 & N5856 );
	assign N6864 = ( N5837 & N3202 );
	assign N6860 = ~( AND3_1815_inw1 | N3202 );
	assign AND4_1809_inw2 = ~( N3202 & N5807 );
	assign N9445 = ~( N3202 & N9093 );
	assign N6203 = ~N3202;
	assign N10415 = ( N3202 | N10290 );
	assign g25_inw1 = ~( N5799 & N3202 );
	assign N9442 = ~( N3628 & N9087 );
	assign N4813 = ~N3628;
	assign AND3_1815_inw1 = ~( N5837 & N5821 );
	assign N6861 = ~( AND3_1816_inw1 | N5837 );
	assign N10289 = ~( AND3_2972_inw1 | N5837 );
	assign AND4_1809_inw1 = ~( N5837 & N5821 );
	assign AND4_1810_inw2 = ~( N5807 & N5837 );
	assign AND4_2971_inw2 = ~( N5821 & N5837 );
	assign N10640 = ~( N5837 & N10563 );
	assign N10915 = ~( N5837 & N10882 );
	assign N10916 = ~( N5837 & N10884 );
	assign N8246 = ~N5837;
	assign g13_inw2 = ~( N5837 & n_322 );
	assign n_328 = ( N5837 & N5821 );
	assign g91_inw1 = ~( N5821 & N5837 );
	assign N6859 = ( N5821 & N3195 );
	assign AND3_1808_inw1 = ~( N5821 & N3195 );
	assign AND4_1805_inw2 = ~( N3195 & N5807 );
	assign N7659 = ( N3195 | N6864 );
	assign OR3_3026_inw1 = ~( N3195 | N6864 );
	assign AND4_1805_inw1 = ~( N5821 & N5799 );
	assign N10639 = ~( N5821 & N10561 );
	assign N11143 = ~( N5821 & N11118 );
	assign N11144 = ~( N5821 & N11120 );
	assign N8245 = ~N5821;
	assign g13_inw1 = ~( N5821 & N5799 );
	assign g79_inw1 = ~( N5821 & N5807 );
	assign N6852 = ( N5807 & N3189 );
	assign N6849 = ~( AND3_1804_inw1 | N3189 );
	assign NOR3_2040_inw1 = ~( N3189 | N6859 );
	assign OR4_2038_inw1 = ~( N3189 | N6859 );
	assign OR4_3025_inw1 = ~( N3189 | N6859 );
	assign AND3_1804_inw1 = ~( N5807 & N5799 );
	assign N6853 = ~( AND3_1808_inw1 | N5807 );
	assign N10638 = ~( N5807 & N10559 );
	assign N11244 = ~( N5807 & N11217 );
	assign N11245 = ~( N5807 & N11219 );
	assign N8244 = ~N5807;
	assign g25_inw2 = ~( N5807 & n_328 );
	assign g91_inw2 = ~( N5807 & N10290 );
	assign N6848 = ( N5799 & N3185 );
	assign NOR4_2041_inw1 = ~( N3185 | N6852 );
	assign n_360 = ( N3185 | N6852 );
	assign N10637 = ~( N5799 & N10557 );
	assign N11027 = ~( N5799 & N10998 );
	assign N11028 = ~( N5799 & N11000 );
	assign N8243 = ~N5799;
	assign g79_inw2 = ~( N5799 & N6866 );
	assign n_325 = ( N3184 | N6848 );
	assign N6865 = ( N5850 & N5789 );
	assign N10710 = ( N5850 & N10589 );
	assign AND3_1798_inw1 = ~( N5850 & N5789 );
	assign AND4_1792_inw1 = ~( N5850 & N5789 );
	assign N10609 = ~( N5850 & N10515 );
	assign N10610 = ~( N5850 & N10517 );
	assign N6761 = ~N5850;
	assign N6844 = ( N5789 & N3178 );
	assign AND3_1797_inw1 = ~( N5789 & N3178 );
	assign AND4_1795_inw2 = ~( N3178 & N5778 );
	assign N8888 = ~( N3178 & N8323 );
	assign N9847 = ~( N3178 & N7650 );
	assign N5943 = ~N3178;
	assign N8887 = ~( N3625 & N8323 );
	assign N9846 = ~( N3625 & N9659 );
	assign N4543 = ~N3625;
	assign AND4_1795_inw1 = ~( N5789 & N5771 );
	assign N8322 = ~( N5789 & N4543 );
	assign N8324 = ~( N5789 & N5943 );
	assign N10845 = ~( N5789 & N10796 );
	assign N10846 = ~( N5789 & N10798 );
	assign N8323 = ~N5789;
	assign N6839 = ( N5778 & N3173 );
	assign N6837 = ~( AND3_1794_inw1 | N3173 );
	assign N8208 = ~( N3173 | N6844 );
	assign OR3_2044_inw1 = ~( N3173 | N6844 );
	assign AND3_1794_inw1 = ~( N5778 & N5771 );
	assign N6840 = ~( AND3_1797_inw1 | N5778 );
	assign N6841 = ~( AND3_1798_inw1 | N5778 );
	assign AND4_1792_inw2 = ~( N5778 & N5771 );
	assign N9273 = ~( N5778 & N8883 );
	assign N9274 = ~( N5778 & N7650 );
	assign N11077 = ~( N5778 & N11040 );
	assign N11078 = ~( N5778 & N11042 );
	assign N8294 = ~N5778;
	assign N6836 = ( N5771 & N3169 );
	assign NOR3_2037_inw1 = ~( N3169 | N6839 );
	assign OR4_2036_inw1 = ~( N3169 | N6839 );
	assign N9271 = ~( N5771 & N8879 );
	assign N9272 = ~( N5771 & N8881 );
	assign N10969 = ~( N5771 & N10934 );
	assign N10970 = ~( N5771 & N10936 );
	assign N8315 = ~N5771;
	assign OR4_2019_inw1 = ~( N3168 | N6836 );
	assign N9318 = ( N8326 & N6957 );
	assign AND3_2117_inw1 = ~( N6957 & N6946 );
	assign N9315 = ~( AND3_2489_inw1 | N6957 );
	assign AND4_2115_inw1 = ~( N6957 & N6946 );
	assign AND4_2475_inw2 = ~( N6946 & N6957 );
	assign AND4_2488_inw2 = ~( N6936 & N6957 );
	assign N10035 = ~( N6957 & N9903 );
	assign N10981 = ~( N6957 & N10953 );
	assign N11031 = ~( N6957 & N11006 );
	assign N9252 = ~N6957;
	assign g17_inw2 = ~( N6957 & n_324 );
	assign n_330 = ( N6957 & N6946 );
	assign g87_inw1 = ~( N6946 & N6957 );
	assign N8355 = ( N4570 & N6946 );
	assign AND3_2114_inw1 = ~( N6946 & N4570 );
	assign AND4_2111_inw2 = ~( N4570 & N6936 );
	assign N8931 = ( N4570 | N8357 );
	assign OR3_2646_inw1 = ~( N4570 | N8357 );
	assign AND3_2489_inw1 = ~( N8326 & N6946 );
	assign AND4_2111_inw1 = ~( N6946 & N6929 );
	assign AND4_2488_inw1 = ~( N8326 & N6946 );
	assign N10034 = ~( N6946 & N9901 );
	assign N11210 = ~( N6946 & N11183 );
	assign N11250 = ~( N6946 & N11231 );
	assign N9251 = ~N6946;
	assign g17_inw1 = ~( N6946 & N6929 );
	assign g83_inw1 = ~( N6946 & N6936 );
	assign N8352 = ( N6936 & N4566 );
	assign N8349 = ~( AND3_2110_inw1 | N4566 );
	assign NOR3_2424_inw1 = ~( N4566 | N8355 );
	assign OR4_2645_inw1 = ~( N4566 | N8355 );
	assign OR4_2667_inw1 = ~( N4566 | N8355 );
	assign AND3_2110_inw1 = ~( N6936 & N6929 );
	assign N8353 = ~( AND3_2114_inw1 | N6936 );
	assign N10033 = ~( N6936 & N9899 );
	assign N11282 = ~( N6936 & N11264 );
	assign N11295 = ~( N6936 & N11290 );
	assign N9250 = ~N6936;
	assign n_324 = ( N6936 & N8326 );
	assign g29_inw2 = ~( N6936 & n_330 );
	assign N8348 = ( N6929 & N4563 );
	assign NOR4_2425_inw1 = ~( N4563 | N8352 );
	assign n_358 = ( N4563 | N8352 );
	assign N10032 = ~( N6929 & N9897 );
	assign N11095 = ~( N6929 & N11065 );
	assign N11145 = ~( N6929 & N11122 );
	assign N9249 = ~N6929;
	assign g83_inw2 = ~( N6929 & N9318 );
	assign n_327 = ( N4562 | N8348 );
	assign N8346 = ( N6923 & N6912 );
	assign N10269 = ( N6923 & N10124 );
	assign AND3_2103_inw1 = ~( N6923 & N6912 );
	assign AND4_2097_inw1 = ~( N6901 & N6923 );
	assign N10748 = ~( N6923 & N10685 );
	assign N10749 = ~( N6923 & N10687 );
	assign N8253 = ~N6923;
	assign N8345 = ( N6912 & N4555 );
	assign AND3_2102_inw1 = ~( N6912 & N4555 );
	assign AND4_2100_inw2 = ~( N4555 & N6901 );
	assign N9570 = ~( N4555 & N9298 );
	assign N10085 = ~( N4555 & N8924 );
	assign N6969 = ~N4555;
	assign N9569 = ~( N4844 & N9298 );
	assign N10084 = ~( N4844 & N9971 );
	assign N5966 = ~N4844;
	assign AND4_2097_inw2 = ~( N6912 & N6894 );
	assign AND4_2100_inw1 = ~( N6912 & N6894 );
	assign N9297 = ~( N6912 & N5966 );
	assign N9299 = ~( N6912 & N6969 );
	assign N10917 = ~( N6912 & N10886 );
	assign N10918 = ~( N6912 & N10888 );
	assign N9298 = ~N6912;
	assign N8340 = ( N6901 & N4549 );
	assign N8338 = ~( AND3_2099_inw1 | N4549 );
	assign N9111 = ~( N4549 | N8345 );
	assign OR3_2420_inw1 = ~( N4549 | N8345 );
	assign AND3_2099_inw1 = ~( N6901 & N6894 );
	assign N8341 = ~( AND3_2102_inw1 | N6901 );
	assign N8342 = ~( AND3_2103_inw1 | N6901 );
	assign N9764 = ~( N6901 & N9565 );
	assign N9765 = ~( N6901 & N8924 );
	assign N11137 = ~( N6901 & N11106 );
	assign N11138 = ~( N6901 & N11108 );
	assign N9294 = ~N6901;
	assign N8337 = ( N6894 & N4545 );
	assign NOR3_2419_inw1 = ~( N4545 | N8340 );
	assign OR4_2418_inw1 = ~( N4545 | N8340 );
	assign N9762 = ~( N6894 & N9561 );
	assign N9763 = ~( N6894 & N9563 );
	assign N11029 = ~( N6894 & N11002 );
	assign N11030 = ~( N6894 & N11004 );
	assign N9290 = ~N6894;
	assign OR4_2371_inw1 = ~( N4544 | N8337 );
	assign N8518 = ( N7180 & N7170 );
	assign N10597 = ( N10381 & N7180 );
	assign AND3_2217_inw1 = ~( N7180 & N7159 );
	assign AND3_3108_inw1 = ~( N10381 & N7180 );
	assign AND4_2211_inw1 = ~( N7180 & N7159 );
	assign AND4_3107_inw1 = ~( N10381 & N7180 );
	assign N10764 = ~( N7180 & N10719 );
	assign N10862 = ~( N7180 & N10823 );
	assign N10863 = ~( N7180 & N10825 );
	assign N9244 = ~N7180;
	assign n_323 = ( N7149 & N7180 );
	assign N8456 = ( N7170 & N4687 );
	assign N8455 = ~( AND3_2179_inw1 | N4687 );
	assign AND4_2177_inw2 = ~( N4687 & N7149 );
	assign N9876 = ~( N4687 & N9721 );
	assign N7573 = ~N4687;
	assign N10668 = ( N4687 | N10597 );
	assign g27_inw1 = ~( N7142 & N4687 );
	assign N9873 = ~( N5030 & N9715 );
	assign N6235 = ~N5030;
	assign AND3_2179_inw1 = ~( N7170 & N7159 );
	assign N8513 = ~( AND3_2217_inw1 | N7170 );
	assign N10596 = ~( AND3_3108_inw1 | N7170 );
	assign AND4_2177_inw1 = ~( N7170 & N7159 );
	assign AND4_2211_inw2 = ~( N7149 & N7170 );
	assign AND4_3107_inw2 = ~( N7159 & N7170 );
	assign N10835 = ~( N7170 & N10775 );
	assign N10986 = ~( N7170 & N10961 );
	assign N10987 = ~( N7170 & N10963 );
	assign N9248 = ~N7170;
	assign g15_inw2 = ~( N7170 & n_323 );
	assign n_329 = ( N7170 & N7159 );
	assign g99_inw1 = ~( N7159 & N7170 );
	assign N8454 = ( N4682 & N7159 );
	assign AND3_2176_inw1 = ~( N7159 & N4682 );
	assign AND4_2173_inw2 = ~( N4682 & N7149 );
	assign N9005 = ( N4682 | N8456 );
	assign OR3_3136_inw1 = ~( N4682 | N8456 );
	assign AND4_2173_inw1 = ~( N7159 & N7142 );
	assign N10834 = ~( N7159 & N10773 );
	assign N11211 = ~( N7159 & N11185 );
	assign N11212 = ~( N7159 & N11187 );
	assign N9247 = ~N7159;
	assign g15_inw1 = ~( N7159 & N7142 );
	assign g81_inw1 = ~( N7159 & N7149 );
	assign N8451 = ( N7149 & N4678 );
	assign N8448 = ~( AND3_2172_inw1 | N4678 );
	assign NOR3_2440_inw1 = ~( N4678 | N8454 );
	assign OR4_2438_inw1 = ~( N4678 | N8454 );
	assign OR4_3135_inw1 = ~( N4678 | N8454 );
	assign AND3_2172_inw1 = ~( N7149 & N7142 );
	assign N8452 = ~( AND3_2176_inw1 | N7149 );
	assign N10833 = ~( N7149 & N10771 );
	assign N11284 = ~( N7149 & N11267 );
	assign N11285 = ~( N7149 & N11269 );
	assign N9246 = ~N7149;
	assign g27_inw2 = ~( N7149 & n_329 );
	assign g99_inw2 = ~( N7149 & N10597 );
	assign N8447 = ( N7142 & N4675 );
	assign NOR4_2441_inw1 = ~( N4675 | N8451 );
	assign n_364 = ( N4675 | N8451 );
	assign N10832 = ~( N7142 & N10769 );
	assign N11098 = ~( N7142 & N11073 );
	assign N11099 = ~( N7142 & N11075 );
	assign N9245 = ~N7142;
	assign g81_inw2 = ~( N7142 & N8518 );
	assign n_326 = ( N4674 | N8447 );
	assign N8442 = ( N7136 & N7125 );
	assign N10867 = ( N7136 & N10784 );
	assign AND3_2164_inw1 = ~( N7136 & N7125 );
	assign AND4_2158_inw1 = ~( N7114 & N7136 );
	assign N10753 = ~( N7136 & N10694 );
	assign N10754 = ~( N7136 & N10696 );
	assign N8252 = ~N7136;
	assign N8441 = ( N7125 & N4667 );
	assign AND3_2163_inw1 = ~( N7125 & N4667 );
	assign AND4_2161_inw2 = ~( N4667 & N7114 );
	assign N9601 = ~( N4667 & N9360 );
	assign N10094 = ~( N4667 & N8996 );
	assign N7187 = ~N4667;
	assign N9600 = ~( N4940 & N9360 );
	assign N10093 = ~( N4940 & N9995 );
	assign N6078 = ~N4940;
	assign AND4_2158_inw2 = ~( N7125 & N7107 );
	assign AND4_2161_inw1 = ~( N7125 & N7107 );
	assign N9359 = ~( N7125 & N6078 );
	assign N9361 = ~( N7125 & N7187 );
	assign N10922 = ~( N7125 & N10895 );
	assign N10923 = ~( N7125 & N10897 );
	assign N9360 = ~N7125;
	assign N8436 = ( N7114 & N4661 );
	assign N8434 = ~( AND3_2160_inw1 | N4661 );
	assign N9173 = ~( N4661 | N8441 );
	assign OR3_2430_inw1 = ~( N4661 | N8441 );
	assign AND3_2160_inw1 = ~( N7114 & N7107 );
	assign N8437 = ~( AND3_2163_inw1 | N7114 );
	assign N8438 = ~( AND3_2164_inw1 | N7114 );
	assign N9797 = ~( N7114 & N9596 );
	assign N9798 = ~( N7114 & N8996 );
	assign N11139 = ~( N7114 & N11110 );
	assign N11140 = ~( N7114 & N11112 );
	assign N9356 = ~N7114;
	assign N8433 = ( N7107 & N4657 );
	assign NOR3_2429_inw1 = ~( N4657 | N8436 );
	assign OR4_2428_inw1 = ~( N4657 | N8436 );
	assign N9795 = ~( N7107 & N9592 );
	assign N9796 = ~( N7107 & N9594 );
	assign N11034 = ~( N7107 & N11011 );
	assign N11035 = ~( N7107 & N11013 );
	assign N9352 = ~N7107;
	assign OR4_2382_inw1 = ~( N4656 | N8433 );
	assign N9904 = ~( N9635 & N9252 );
	assign N9903 = ~N9635;
	assign N9285 = ~( g87_inw1 | g87_inw2 );
	assign N10105 = ( N9925 & N9894 );
	assign N10106 = ( N9925 & N9895 );
	assign N10107 = ( N9925 & N9896 );
	assign N10108 = ( N9925 & N8253 );
	assign N10130 = ( N9768 & N9925 );
	assign N10124 = ~N9925;
	assign N11336 = ~( N11323 & N11283 );
	assign N11337 = ~N11323;
	assign N9632 = ~( OR3_2646_inw1 & N9287 );
	assign N10119 = ~( OR3_2893_inw1 & N10043 );
	assign N10148 = ~( OR3_2907_inw1 & N10061 );
	assign N11252 = ~( OR4_3452_inw1 & OR4_3452_inw2 );
	assign OR4_2645_inw2 = ~( N8356 | N9286 );
	assign OR4_2892_inw2 = ~( N10040 | N10041 );
	assign OR4_2906_inw2 = ~( N10058 | N10059 );
	assign N10133 = ( N9932 & N8898 );
	assign N10131 = ~N9932;
	assign OR4_3452_inw1 = ~( N11222 | N11223 );
	assign N10015 = ~( g5_inw1 | g5_inw2 );
	assign N10022 = ~( g75_inw1 | g75_inw2 );
	assign N1489 = N1113;
	assign AND4_1887_inw2 = ~( N3373 & N6047 );
	assign N5751 = ~( N5185 & N5186 );
	assign N6056 = ~( N5320 & N5321 );
	assign N6052 = ~( N5318 & N5319 );
	assign N7104 = ~( g40_inw1 | g40_inw2 );
	assign N7103 = ( N6041 & N3371 );
	assign N5755 = ~( N5187 & N5188 );
	assign N6047 = ~( N5316 & N5317 );
	assign n_334 = ( N3370 | N7103 );
	assign N6041 = ~( N5314 & N5315 );
	assign n_342 = ( N3365 | N7064 );
	assign N6003 = ~( N5289 & N5290 );
	assign N6145 = ~( N5432 & N5433 );
	assign AND4_1869_inw2 = ~( N3364 & N5996 );
	assign N6021 = ~( N5297 & N5298 );
	assign N6252 = ~( N5584 & N5585 );
	assign N6000 = ~( N5287 & N5288 );
	assign N7061 = ~( g44_inw1 | g44_inw2 );
	assign N7060 = ( N5991 & N3362 );
	assign N5996 = ~( N5285 & N5286 );
	assign N6249 = ~( N5586 & N5587 );
	assign OR4_2027_inw1 = ~( N3361 | N7060 );
	assign N5991 = ~( N5283 & N5284 );
	assign N5766 = ~( N5192 & N5193 );
	assign N6199 = ~( N5474 & N5475 );
	assign N6196 = ~( N5476 & N5477 );
	assign N5740 = ~( N5180 & N5181 );
	assign N5744 = ~( N5182 & N5183 );
	assign N4803 = ~( N4326 & N4327 );
	assign N4806 = ~( N4333 & N4334 );
	assign AND3_2075_inw1 = ~( N5740 & N5736 );
	assign AND3_2353_inw1 = ~( N5736 & N6800 );
	assign N6797 = ~N5736;
	assign AND3_2077_inw1 = ~( N5751 & N5747 );
	assign AND3_2355_inw1 = ~( N5747 & N6806 );
	assign N6803 = ~N5747;
	assign n_339 = ( N6059 & N6056 );
	assign g36_inw2 = ~( N7106 | n_334 );
	assign N6137 = ~( N5429 & N4751 );
	assign N6022 = ~( N5299 & N5300 );
	assign N7067 = ~( g62_inw1 | g62_inw2 );
	assign AND4_1873_inw2 = ~( N3368 & N6009 );
	assign N6018 = ~( N5295 & N5296 );
	assign N6141 = ~( N5430 & N5431 );
	assign N6014 = ~( N5293 & N5294 );
	assign N7065 = ~( g59_inw1 | g59_inw2 );
	assign N7064 = ( N6003 & N3366 );
	assign N6009 = ~( N5291 & N5292 );
	assign N5758 = ~( N5189 & N4502 );
	assign N5762 = ~( N5190 & N5191 );
	assign N6079 = ~( N5363 & N4694 );
	assign g43_inw2 = ~( n_337 & n_338 );
	assign N6083 = ~( N5364 & N5365 );
	assign N6087 = ~( N5366 & N5367 );
	assign N4997 = ~( N4411 & N4412 );
	assign N6166 = ~( N5451 & N4776 );
	assign g62_inw2 = ~( n_336 & n_346 );
	assign N6170 = ~( N5452 & N5453 );
	assign N6174 = ~( N5454 & N5455 );
	assign N6266 = ~( N5602 & N5603 );
	assign N6263 = ~( N5604 & N5605 );
	assign N6127 = ~( N5425 & N4746 );
	assign AND4_2240_inw2 = ~( N4766 & N7364 );
	assign N6131 = ~( N5426 & N5427 );
	assign N7373 = ~( N6687 & N6161 );
	assign N7369 = ~( N6686 & N6159 );
	assign N8552 = ~( g67_inw1 | g67_inw2 );
	assign N8551 = ( N7358 & N4762 );
	assign N7331 = ~( N6668 & N6136 );
	assign N7364 = ~( N6685 & N6157 );
	assign n_343 = ( N4637 | N8415 );
	assign N7080 = ~( N6597 & N6030 );
	assign N7322 = ~( N6125 & N6661 );
	assign AND4_2151_inw2 = ~( N4635 & N7073 );
	assign N6246 = ~( N5571 & N5572 );
	assign N7098 = ~( N6604 & N6038 );
	assign N7077 = ~( N6596 & N6028 );
	assign N8410 = ~( g53_inw1 | g53_inw2 );
	assign N8409 = ( N7068 & N4632 );
	assign N6243 = ~( N5573 & N5574 );
	assign N7073 = ~( N6595 & N6026 );
	assign OR4_2378_inw1 = ~( N4630 | N8409 );
	assign N7068 = ~( N6594 & N6024 );
	assign n_344 = ( N4760 | N8551 );
	assign N7358 = ~( N6683 & N6684 );
	assign AND4_2236_inw2 = ~( N4759 & N7351 );
	assign N7376 = ~( N6688 & N6689 );
	assign N7577 = ~( N6741 & N6742 );
	assign N7355 = ~( N6681 & N6682 );
	assign N8546 = ~( g56_inw1 | g56_inw2 );
	assign N8545 = ( N7346 & N4757 );
	assign N7351 = ~( N6679 & N6680 );
	assign N7574 = ~( N6743 & N6744 );
	assign OR4_2392_inw1 = ~( N4756 | N8545 );
	assign N7346 = ~( N6677 & N6678 );
	assign N7213 = ~( N6647 & N6648 );
	assign N7569 = ~( N6733 & N6734 );
	assign N7566 = ~( N6735 & N6736 );
	assign N7314 = ~( N6658 & N6122 );
	assign N7099 = ~( N6605 & N6606 );
	assign N8418 = ~( g66_inw1 | g66_inw2 );
	assign AND4_2155_inw2 = ~( N4640 & N7086 );
	assign N7095 = ~( N6602 & N6603 );
	assign N7318 = ~( N6659 & N6660 );
	assign N7091 = ~( N6600 & N6601 );
	assign N8416 = ~( g63_inw1 | g63_inw2 );
	assign N8415 = ( N7080 & N4638 );
	assign N7086 = ~( N6598 & N6599 );
	assign N7194 = ~( N6639 & N6091 );
	assign N7198 = ~( N6640 & N6641 );
	assign N7202 = ~( N6642 & N6643 );
	assign N7205 = ~( N6644 & N6097 );
	assign N7209 = ~( N6645 & N6646 );
	assign N7563 = ~( N6729 & N6730 );
	assign N7560 = ~( N6731 & N6732 );
	assign N7394 = ~( N6706 & N6186 );
	assign g66_inw2 = ~( n_347 & n_348 );
	assign N7398 = ~( N6707 & N6708 );
	assign N7402 = ~( N6709 & N6710 );
	assign N7591 = ~( N6755 & N6756 );
	assign N7588 = ~( N6757 & N6758 );
	assign N6177 = ~( N5456 & N5457 );
	assign N7387 = ~( N6702 & N6703 );
	assign N7391 = ~( N6704 & N6705 );
	assign N7585 = ~( N6751 & N6752 );
	assign N7582 = ~( N6753 & N6754 );
	assign N8554 = ~( g70_inw1 | g70_inw2 );
	assign NOR3_2424_invw = ~( NOR3_2424_inw1 & N8356 );
	assign OR4_2667_inw2 = ~( N8356 | N9315 );
	assign N8354 = ~( AND4_2115_inw1 | AND4_2115_inw2 );
	assign N9979 = ~( N9691 & N9863 );
	assign N9691 = ~( N9146 & N8717 );
	assign N8351 = ~( g29_inw1 | g29_inw2 );
	assign N10857 = ~( N8326 & N10815 );
	assign N10919 = ~( N8326 & N10890 );
	assign N9741 = ~N8326;
	assign N10192 = ~( N9976 & N10086 );
	assign N9976 = ~( N9679 & N7552 );
	assign n_341 = ( N7377 & N7373 );
	assign N10549 = ( N5165 & N10367 );
	assign N10631 = ( N5165 & N10550 );
	assign N9429 = ~( N9065 & N8610 );
	assign N10551 = ( N10354 & N3126 );
	assign N10705 = ( N3126 & N10583 );
	assign N8610 = ~( N7444 & N3126 );
	assign N4784 = ( N3126 | N3122 );
	assign n_316 = ( N3126 | N8818 );
	assign N9064 = ~( N4303 & N8607 );
	assign N5469 = ~N4303;
	assign N10730 = ( N5178 & N10583 );
	assign N8609 = ~N7444;
	assign N10628 = ( N10546 | N10451 );
	assign N5631 = ~( N5324 & N4653 );
	assign g32_inw2 = ~( n_331 | n_332 );
	assign N8262 = ( N3122 & N6762 );
	assign N8269 = ( N3122 & N6784 );
	assign N8818 = ( N7609 & N3122 );
	assign N4473 = ~N3122;
	assign N10357 = ~( N10271 & N10212 );
	assign N10360 = ~( N10272 & N10213 );
	assign N10212 = ~( N10070 & N3954 );
	assign N10213 = ~( N10073 & N3954 );
	assign N10839 = ( N10731 | N10588 );
	assign N10070 = ~( N9955 & N9836 );
	assign N10073 = ~( N9956 & N9838 );
	assign N10588 = ( N10367 & N3135 );
	assign N9836 = ~( N9426 & N3135 );
	assign N9838 = ~( N9429 & N3135 );
	assign N8421 = ( N3375 & N7100 );
	assign N8960 = ( N3375 & N7852 );
	assign N4653 = ~N3375;
	assign N5735 = ~N5177;
	assign N8608 = ~( N7441 & N5469 );
	assign N8607 = ~N7441;
	assign N10140 = ~( OR4_2905_inw1 & OR4_2905_inw2 );
	assign N10233 = ( N10139 | N10054 );
	assign N10139 = ( N9785 & N10053 );
	assign g32_inw1 = ~( N10017 | N9734 );
	assign N6768 = ~( AND4_1753_inw1 | AND4_1753_inw2 );
	assign N6772 = ~( AND4_1757_inw1 | AND4_1757_inw2 );
	assign N6773 = ~( AND4_1758_inw1 | AND4_1758_inw2 );
	assign N10279 = ~( AND4_2965_inw1 | AND4_2965_inw2 );
	assign N10717 = ~( N10644 & N10571 );
	assign N11168 = ~( N11141 & N11115 );
	assign N11171 = ~( N11142 & N11117 );
	assign N10571 = ~( N10425 & N8250 );
	assign N11115 = ~( N11044 & N8250 );
	assign N11117 = ~( N11047 & N8250 );
	assign N6784 = ~( g11_inw1 | g11_inw2 );
	assign N6762 = ~( g77_inw1 | g77_inw2 );
	assign N10278 = ~( g95_inw1 | g95_inw2 );
	assign g7_inw1 = ~( N6767 | N6768 );
	assign NOR3_2032_invw = ~( NOR3_2032_inw1 & N6778 );
	assign N8114 = ~( OR4_2030_inw1 & OR4_2030_inw2 );
	assign N10422 = ~( OR4_3029_inw1 & OR4_3029_inw2 );
	assign AND3_3130_inw1 = ~( N886 & N887 );
	assign N9068 = ( N7613 | N6783 );
	assign N10641 = ~( N10565 & N10466 );
	assign N10789 = ~( N10737 & N10672 );
	assign N10792 = ~( N10738 & N10674 );
	assign N10466 = ~( N10141 & N8247 );
	assign N10672 = ~( N10509 & N8247 );
	assign N10674 = ~( N10512 & N8247 );
	assign OR4_2030_inw2 = ~( N6778 | N6779 );
	assign OR4_3029_inw2 = ~( N6778 | N10279 );
	assign N9646 = ~( N9073 & N9435 );
	assign N9073 = ~( N8131 & N6195 );
	assign N10573 = ~( N10428 & N8251 );
	assign N10572 = ~N10428;
	assign N6769 = ~( g9_inw1 | g9_inw2 );
	assign N9642 = ~( N9067 & N9432 );
	assign N9067 = ~( N8114 & N4795 );
	assign N10425 = ~( OR3_3030_inw1 & N10280 );
	assign N10718 = ~( N10645 & N10573 );
	assign N10928 = ~( N10909 & N10873 );
	assign N10931 = ~( N10910 & N10875 );
	assign N10873 = ~( N10789 & N8251 );
	assign N10875 = ~( N10792 & N8251 );
	assign N9960 = ~( N9646 & N7613 );
	assign N9074 = ~N7613;
	assign NOR4_2033_inw2 = ~( N6771 | N6772 );
	assign g93_inw1 = ~( N6771 | N6772 );
	assign g103_inw1 = ~( N6771 | N6772 );
	assign N10716 = ~( N10643 & N10569 );
	assign N11260 = ~( N11242 & N11214 );
	assign N11261 = ~( N11243 & N11216 );
	assign N10569 = ~( N10422 & N8249 );
	assign N11214 = ~( N11168 & N8249 );
	assign N11216 = ~( N11171 & N8249 );
	assign NOR4_2033_invw = ~( NOR4_2033_inw1 & NOR4_2033_inw2 );
	assign g93_inw2 = ~( N10278 | n_362 );
	assign g103_inw2 = ~( N6773 | n_362 );
	assign N10715 = ~( N10642 & N10567 );
	assign N11044 = ~( N11023 & N10989 );
	assign N11047 = ~( N11024 & N10991 );
	assign N10567 = ~( N10419 & N8248 );
	assign N10989 = ~( N10928 & N8248 );
	assign N10991 = ~( N10931 & N8248 );
	assign g7_inw2 = ~( N6769 | n_319 );
	assign N9089 = ( N7659 | N6866 );
	assign N6855 = ~( AND4_1810_inw1 | AND4_1810_inw2 );
	assign N10288 = ~( AND4_2971_inw1 | AND4_2971_inw2 );
	assign N10632 = ~( N10552 & N10456 );
	assign N10800 = ~( N10746 & N10682 );
	assign N10803 = ~( N10747 & N10684 );
	assign N10456 = ~( N10148 & N8242 );
	assign N10682 = ~( N10519 & N8242 );
	assign N10684 = ~( N10522 & N8242 );
	assign NOR3_2040_invw = ~( NOR3_2040_inw1 & N6860 );
	assign OR4_2038_inw2 = ~( N6860 | N6861 );
	assign OR4_3025_inw2 = ~( N6860 | N10288 );
	assign N6854 = ~( AND4_1809_inw1 | AND4_1809_inw2 );
	assign N9667 = ~( N9094 & N9445 );
	assign N9094 = ~( N8183 & N6203 );
	assign N10564 = ~( N10415 & N8246 );
	assign N10563 = ~N10415;
	assign N6851 = ~( g25_inw1 | g25_inw2 );
	assign N9663 = ~( N9088 & N9442 );
	assign N9088 = ~( N8166 & N4813 );
	assign N10412 = ~( OR3_3026_inw1 & N10289 );
	assign N10714 = ~( N10640 & N10564 );
	assign N10938 = ~( N10915 & N10883 );
	assign N10941 = ~( N10916 & N10885 );
	assign N10883 = ~( N10800 & N8246 );
	assign N10885 = ~( N10803 & N8246 );
	assign N6881 = ~( g13_inw1 | g13_inw2 );
	assign N10287 = ~( g91_inw1 | g91_inw2 );
	assign N6850 = ~( AND4_1805_inw1 | AND4_1805_inw2 );
	assign N9970 = ~( N9667 & N7659 );
	assign N9095 = ~N7659;
	assign N10713 = ~( N10639 & N10562 );
	assign N11174 = ~( N11143 & N11119 );
	assign N11177 = ~( N11144 & N11121 );
	assign N10562 = ~( N10412 & N8245 );
	assign N11119 = ~( N11050 & N8245 );
	assign N11121 = ~( N11053 & N8245 );
	assign N6845 = ~( g79_inw1 | g79_inw2 );
	assign g19_inw1 = ~( N6849 | N6850 );
	assign N8166 = ~( OR4_2038_inw1 & OR4_2038_inw2 );
	assign N10409 = ~( OR4_3025_inw1 & OR4_3025_inw2 );
	assign NOR4_2041_inw2 = ~( N6853 | N6854 );
	assign g89_inw1 = ~( N6853 | N6854 );
	assign g101_inw1 = ~( N6853 | N6854 );
	assign N10712 = ~( N10638 & N10560 );
	assign N11262 = ~( N11244 & N11218 );
	assign N11263 = ~( N11245 & N11220 );
	assign N10560 = ~( N10409 & N8244 );
	assign N11218 = ~( N11174 & N8244 );
	assign N11220 = ~( N11177 & N8244 );
	assign NOR4_2041_invw = ~( NOR4_2041_inw1 & NOR4_2041_inw2 );
	assign g89_inw2 = ~( N10287 | n_360 );
	assign g101_inw2 = ~( N6855 | n_360 );
	assign N10711 = ~( N10637 & N10558 );
	assign N11050 = ~( N11027 & N10999 );
	assign N11053 = ~( N11028 & N11001 );
	assign N10558 = ~( N10406 & N8243 );
	assign N10999 = ~( N10938 & N8243 );
	assign N11001 = ~( N10941 & N8243 );
	assign g19_inw2 = ~( N6851 | n_325 );
	assign N9079 = ( N7650 | N6865 );
	assign N8204 = ~( OR3_2044_inw1 & N6865 );
	assign N10763 = ( N10710 | N10556 );
	assign N6833 = ~( AND4_1792_inw1 | AND4_1792_inw2 );
	assign N10675 = ~( N10609 & N10516 );
	assign N10678 = ~( N10610 & N10518 );
	assign N10556 = ( N10375 & N6761 );
	assign N10516 = ~( N10318 & N6761 );
	assign N10518 = ~( N10321 & N6761 );
	assign N6838 = ~( AND4_1795_inw1 | AND4_1795_inw2 );
	assign N9243 = ~( N8324 & N8888 );
	assign N9964 = ~( N9662 & N9847 );
	assign N9662 = ~( N8208 & N5943 );
	assign N9275 = ~( N8322 & N8887 );
	assign N9961 = ~( N9660 & N9846 );
	assign N9660 = ~( N9079 & N4543 );
	assign N10876 = ~( N10845 & N10797 );
	assign N10879 = ~( N10846 & N10799 );
	assign N10797 = ~( N10675 & N8323 );
	assign N10799 = ~( N10678 & N8323 );
	assign OR4_2019_inw2 = ~( N6837 | N6838 );
	assign N8886 = ~( N8208 & N8294 );
	assign N7650 = ~N8208;
	assign NOR3_2037_invw = ~( NOR3_2037_inw1 & N6840 );
	assign OR4_2036_inw2 = ~( N6840 | N6841 );
	assign N9540 = ~( N9273 & N8884 );
	assign N9556 = ~( N9274 & N8886 );
	assign N11100 = ~( N11077 & N11041 );
	assign N11103 = ~( N11078 & N11043 );
	assign N8884 = ~( N8204 & N8294 );
	assign N11041 = ~( N10992 & N8294 );
	assign N11043 = ~( N10995 & N8294 );
	assign N8146 = ~( OR4_2036_inw1 & OR4_2036_inw2 );
	assign N9539 = ~( N9271 & N8880 );
	assign N9555 = ~( N9272 & N8882 );
	assign N10992 = ~( N10969 & N10935 );
	assign N10995 = ~( N10970 & N10937 );
	assign N8880 = ~( N8146 & N8315 );
	assign N8882 = ~( N8156 & N8315 );
	assign N10935 = ~( N10876 & N8315 );
	assign N10937 = ~( N10879 & N8315 );
	assign N7649 = ~( OR4_2019_inw1 & OR4_2019_inw2 );
	assign N9682 = ( N8931 | N9318 );
	assign N9314 = ~( AND4_2488_inw1 | AND4_2488_inw2 );
	assign N10112 = ~( N10035 & N9904 );
	assign N11008 = ~( N10981 & N10954 );
	assign N11062 = ~( N11031 & N11007 );
	assign N10954 = ~( N10892 & N9252 );
	assign N11007 = ~( N10950 & N9252 );
	assign N9280 = ~( g17_inw1 | g17_inw2 );
	assign N8350 = ~( AND4_2111_inw1 | AND4_2111_inw2 );
	assign N10196 = ~( N9979 & N8931 );
	assign N9692 = ~N8931;
	assign N10111 = ~( N10034 & N9902 );
	assign N11233 = ~( N11210 & N11184 );
	assign N11272 = ~( N11250 & N11232 );
	assign N9902 = ~( N9632 & N9251 );
	assign N11184 = ~( N11124 & N9251 );
	assign N11232 = ~( N11180 & N9251 );
	assign N9307 = ~( g83_inw1 | g83_inw2 );
	assign g23_inw1 = ~( N8349 | N8350 );
	assign N9629 = ~( OR4_2645_inw1 & OR4_2645_inw2 );
	assign N9679 = ~( OR4_2667_inw1 & OR4_2667_inw2 );
	assign NOR4_2425_inw2 = ~( N8353 | N8354 );
	assign g85_inw1 = ~( N8353 | N8354 );
	assign g107_inw1 = ~( N8353 | N8354 );
	assign N10110 = ~( N10033 & N9900 );
	assign N11292 = ~( N11282 & N11265 );
	assign N11307 = ~( N11295 & N11291 );
	assign N9900 = ~( N9629 & N9250 );
	assign N11265 = ~( N11233 & N9250 );
	assign N11291 = ~( N11272 & N9250 );
	assign NOR4_2425_invw = ~( NOR4_2425_inw1 & NOR4_2425_inw2 );
	assign g85_inw2 = ~( N9285 | n_358 );
	assign g107_inw2 = ~( N9314 | n_358 );
	assign N10109 = ~( N10032 & N9898 );
	assign N11124 = ~( N11095 & N11066 );
	assign N11180 = ~( N11145 & N11123 );
	assign N9898 = ~( N9626 & N9249 );
	assign N11066 = ~( N11008 & N9249 );
	assign N11123 = ~( N11062 & N9249 );
	assign g23_inw2 = ~( N8351 | n_327 );
	assign N9671 = ( N8924 | N8346 );
	assign N9107 = ~( OR3_2420_inw1 & N8346 );
	assign N10353 = ( N10269 | N10108 );
	assign N8333 = ~( AND4_2097_inw1 | AND4_2097_inw2 );
	assign N10806 = ~( N10748 & N10686 );
	assign N10809 = ~( N10749 & N10688 );
	assign N10686 = ~( N10525 & N8253 );
	assign N10688 = ~( N10528 & N8253 );
	assign N8339 = ~( AND4_2100_inw1 | AND4_2100_inw2 );
	assign N9742 = ~( N9299 & N9570 );
	assign N10189 = ~( N9974 & N10085 );
	assign N9974 = ~( N9111 & N6969 );
	assign N9766 = ~( N9297 & N9569 );
	assign N10186 = ~( N9972 & N10084 );
	assign N9972 = ~( N9671 & N5966 );
	assign N10944 = ~( N10917 & N10887 );
	assign N10947 = ~( N10918 & N10889 );
	assign N10887 = ~( N10806 & N9298 );
	assign N10889 = ~( N10809 & N9298 );
	assign OR4_2371_inw2 = ~( N8338 | N8339 );
	assign N9568 = ~( N9111 & N9294 );
	assign N8924 = ~N9111;
	assign NOR3_2419_invw = ~( NOR3_2419_inw1 & N8341 );
	assign OR4_2418_inw2 = ~( N8341 | N8342 );
	assign N9895 = ~( N9764 & N9566 );
	assign N9924 = ~( N9765 & N9568 );
	assign N11156 = ~( N11137 & N11107 );
	assign N11159 = ~( N11138 & N11109 );
	assign N9566 = ~( N9107 & N9294 );
	assign N11107 = ~( N11056 & N9294 );
	assign N11109 = ~( N11059 & N9294 );
	assign N9099 = ~( OR4_2418_inw1 & OR4_2418_inw2 );
	assign N9894 = ~( N9762 & N9562 );
	assign N9923 = ~( N9763 & N9564 );
	assign N11056 = ~( N11029 & N11003 );
	assign N11059 = ~( N11030 & N11005 );
	assign N9562 = ~( N9099 & N9290 );
	assign N9564 = ~( N9103 & N9290 );
	assign N11003 = ~( N10944 & N9290 );
	assign N11005 = ~( N10947 & N9290 );
	assign N8898 = ~( OR4_2371_inw1 & OR4_2371_inw2 );
	assign N9717 = ( N9005 | N8518 );
	assign N8507 = ~( AND4_2211_inw1 | AND4_2211_inw2 );
	assign N10595 = ~( AND4_3107_inw1 | AND4_3107_inw2 );
	assign N10827 = ~( N10764 & N10720 );
	assign N10899 = ~( N10862 & N10824 );
	assign N10902 = ~( N10863 & N10826 );
	assign N10720 = ~( N10381 & N9244 );
	assign N10824 = ~( N10698 & N9244 );
	assign N10826 = ~( N10701 & N9244 );
	assign NOR3_2440_invw = ~( NOR3_2440_inw1 & N8455 );
	assign OR4_2438_inw2 = ~( N8455 | N8513 );
	assign OR4_3135_inw2 = ~( N8455 | N10595 );
	assign N8453 = ~( AND4_2177_inw1 | AND4_2177_inw2 );
	assign N10003 = ~( N9722 & N9876 );
	assign N9722 = ~( N9220 & N7573 );
	assign N10776 = ~( N10668 & N9248 );
	assign N10775 = ~N10668;
	assign N8450 = ~( g27_inw1 | g27_inw2 );
	assign N9999 = ~( N9716 & N9873 );
	assign N9716 = ~( N9203 & N6235 );
	assign N10665 = ~( OR3_3136_inw1 & N10596 );
	assign N10871 = ~( N10835 & N10776 );
	assign N11015 = ~( N10986 & N10962 );
	assign N11018 = ~( N10987 & N10964 );
	assign N10962 = ~( N10899 & N9248 );
	assign N10964 = ~( N10902 & N9248 );
	assign N8444 = ~( g15_inw1 | g15_inw2 );
	assign N10594 = ~( g99_inw1 | g99_inw2 );
	assign N8449 = ~( AND4_2173_inw1 | AND4_2173_inw2 );
	assign N10206 = ~( N10003 & N9005 );
	assign N9723 = ~N9005;
	assign N10870 = ~( N10834 & N10774 );
	assign N11236 = ~( N11211 & N11186 );
	assign N11239 = ~( N11212 & N11188 );
	assign N10774 = ~( N10665 & N9247 );
	assign N11186 = ~( N11127 & N9247 );
	assign N11188 = ~( N11130 & N9247 );
	assign N8497 = ~( g81_inw1 | g81_inw2 );
	assign g21_inw1 = ~( N8448 | N8449 );
	assign N9203 = ~( OR4_2438_inw1 & OR4_2438_inw2 );
	assign N10662 = ~( OR4_3135_inw1 & OR4_3135_inw2 );
	assign NOR4_2441_inw2 = ~( N8452 | N8453 );
	assign g97_inw1 = ~( N8452 | N8453 );
	assign g105_inw1 = ~( N8452 | N8453 );
	assign N10869 = ~( N10833 & N10772 );
	assign N11293 = ~( N11284 & N11268 );
	assign N11294 = ~( N11285 & N11270 );
	assign N10772 = ~( N10662 & N9246 );
	assign N11268 = ~( N11236 & N9246 );
	assign N11270 = ~( N11239 & N9246 );
	assign NOR4_2441_invw = ~( NOR4_2441_inw1 & NOR4_2441_inw2 );
	assign g97_inw2 = ~( N10594 | n_364 );
	assign g105_inw2 = ~( N8507 | n_364 );
	assign N10868 = ~( N10832 & N10770 );
	assign N11127 = ~( N11098 & N11074 );
	assign N11130 = ~( N11099 & N11076 );
	assign N10770 = ~( N10659 & N9245 );
	assign N11074 = ~( N11015 & N9245 );
	assign N11076 = ~( N11018 & N9245 );
	assign g21_inw2 = ~( N8450 | n_326 );
	assign N9707 = ( N8996 | N8442 );
	assign N9169 = ~( OR3_2430_inw1 & N8442 );
	assign N10908 = ( N10867 | N10768 );
	assign N8430 = ~( AND4_2158_inw1 | AND4_2158_inw2 );
	assign N10817 = ~( N10753 & N10695 );
	assign N10820 = ~( N10754 & N10697 );
	assign N10768 = ( N10652 & N8252 );
	assign N10695 = ~( N10536 & N8252 );
	assign N10697 = ~( N10539 & N8252 );
	assign N8435 = ~( AND4_2161_inw1 | AND4_2161_inw2 );
	assign N9739 = ~( N9361 & N9601 );
	assign N10200 = ~( N9998 & N10094 );
	assign N9998 = ~( N9173 & N7187 );
	assign N9799 = ~( N9359 & N9600 );
	assign N10197 = ~( N9996 & N10093 );
	assign N9996 = ~( N9707 & N6078 );
	assign N10955 = ~( N10922 & N10896 );
	assign N10958 = ~( N10923 & N10898 );
	assign N10896 = ~( N10817 & N9360 );
	assign N10898 = ~( N10820 & N9360 );
	assign OR4_2382_inw2 = ~( N8434 | N8435 );
	assign N9599 = ~( N9173 & N9356 );
	assign N8996 = ~N9173;
	assign NOR3_2429_invw = ~( NOR3_2429_inw1 & N8437 );
	assign OR4_2428_inw2 = ~( N8437 | N8438 );
	assign N9891 = ~( N9797 & N9597 );
	assign N9946 = ~( N9798 & N9599 );
	assign N11162 = ~( N11139 & N11111 );
	assign N11165 = ~( N11140 & N11113 );
	assign N9597 = ~( N9169 & N9356 );
	assign N11111 = ~( N11067 & N9356 );
	assign N11113 = ~( N11070 & N9356 );
	assign N9161 = ~( OR4_2428_inw1 & OR4_2428_inw2 );
	assign N9890 = ~( N9795 & N9593 );
	assign N9945 = ~( N9796 & N9595 );
	assign N11067 = ~( N11034 & N11012 );
	assign N11070 = ~( N11035 & N11014 );
	assign N9593 = ~( N9161 & N9352 );
	assign N9595 = ~( N9165 & N9352 );
	assign N11012 = ~( N10955 & N9352 );
	assign N11014 = ~( N10958 & N9352 );
	assign N8963 = ~( OR4_2382_inw1 & OR4_2382_inw2 );
	assign N10350 = ( N10266 | N10105 );
	assign N10351 = ( N10267 | N10106 );
	assign N10352 = ( N10268 | N10107 );
	assign N10381 = ( N10292 | N10130 );
	assign N10266 = ( N10026 & N10124 );
	assign N10267 = ( N10028 & N10124 );
	assign N10268 = ( N9742 & N10124 );
	assign N10292 = ( N8898 & N10124 );
	assign N11341 = ~( N11336 & N11339 );
	assign N11339 = ~( N11252 & N11337 );
	assign N9901 = ~N9632;
	assign N11280 = ( N10119 & N11262 );
	assign N11154 = ~( AND3_3404_inw1 | N10119 );
	assign N11155 = ~( AND3_3405_inw1 | N10119 );
	assign N10283 = ~N10119;
	assign N10291 = ( N6881 & N10148 );
	assign N10455 = ~N10148;
	assign N11283 = ~N11252;
	assign N10116 = ~( OR4_2892_inw1 & OR4_2892_inw2 );
	assign N10141 = ~( OR4_2906_inw1 & OR4_2906_inw2 );
	assign N10301 = ( N10230 | N10133 );
	assign N10230 = ( N9768 & N10131 );
	assign g3_inw1 = ~( N10014 | N10015 );
	assign g73_inw1 = ~( N10021 | N10022 );
	assign N7105 = ~( AND4_1887_inw1 | AND4_1887_inw2 );
	assign AND3_2354_inw1 = ~( N6803 & N5751 );
	assign N6806 = ~N5751;
	assign n_337 = ( N6056 & N6052 );
	assign AND4_1887_inw1 = ~( N6052 & N6041 );
	assign g46_inw1 = ~( N6052 & N6047 );
	assign g36_inw1 = ~( N7104 | N7105 );
	assign N8282 = ~( AND3_2077_inw1 | N5755 );
	assign N8283 = ~( AND3_2078_inw1 | N5755 );
	assign N8276 = ~N5755;
	assign g40_inw1 = ~( N6047 & N6041 );
	assign g46_inw2 = ~( N6041 & n_339 );
	assign g52_inw2 = ~( N7067 | n_342 );
	assign AND4_1873_inw1 = ~( N6014 & N6003 );
	assign g39_inw1 = ~( N6009 & N6003 );
	assign g59_inw1 = ~( N6009 & N6003 );
	assign N8539 = ~( AND3_2231_inw1 | N6145 );
	assign N8540 = ~( AND3_2232_inw1 | N6145 );
	assign N8537 = ~N6145;
	assign N7062 = ~( AND4_1869_inw1 | AND4_1869_inw2 );
	assign AND4_1866_inw1 = ~( N6021 & N6000 );
	assign N8216 = ~( N6252 & N7556 );
	assign N7557 = ~N6252;
	assign AND4_1869_inw1 = ~( N6000 & N5991 );
	assign OR4_2027_inw2 = ~( N7061 | N7062 );
	assign AND4_1866_inw2 = ~( N5996 & N5991 );
	assign g44_inw1 = ~( N5996 & N5991 );
	assign N8217 = ~( N6249 & N7557 );
	assign N7556 = ~N6249;
	assign N7825 = ~( OR4_2027_inw1 & OR4_2027_inw2 );
	assign N8284 = ~( AND3_2079_inw1 | N5766 );
	assign N8285 = ~( AND3_2080_inw1 | N5766 );
	assign N8278 = ~N5766;
	assign N8144 = ~( N6199 & N7477 );
	assign N7478 = ~N6199;
	assign N8145 = ~( N6196 & N7478 );
	assign N7477 = ~N6196;
	assign AND3_2352_inw1 = ~( N6797 & N5740 );
	assign N6800 = ~N5740;
	assign N8280 = ~( AND3_2075_inw1 | N5744 );
	assign N8281 = ~( AND3_2076_inw1 | N5744 );
	assign N8274 = ~N5744;
	assign N10036 = ~( N4803 & N9906 );
	assign N5769 = ~N4803;
	assign N10037 = ~( N4806 & N9908 );
	assign N5770 = ~N4806;
	assign N8862 = ~( AND3_2353_inw1 | N8274 );
	assign AND3_2076_inw1 = ~( N6800 & N6797 );
	assign N8864 = ~( AND3_2355_inw1 | N8276 );
	assign AND3_2078_inw1 = ~( N6806 & N6803 );
	assign N7852 = ~( g36_inw1 & g36_inw2 );
	assign AND3_2231_inw1 = ~( N6141 & N6137 );
	assign AND3_2391_inw1 = ~( N6137 & N7337 );
	assign N7334 = ~N6137;
	assign n_335 = ( N7057 & N6022 );
	assign N7066 = ~( AND4_1873_inw1 | AND4_1873_inw2 );
	assign n_336 = ( N6018 & N6014 );
	assign AND3_2390_inw1 = ~( N7334 & N6141 );
	assign N7337 = ~N6141;
	assign g52_inw1 = ~( N7065 | N7066 );
	assign AND3_2079_inw1 = ~( N5762 & N5758 );
	assign AND3_2357_inw1 = ~( N5758 & N6812 );
	assign N6809 = ~N5758;
	assign AND3_2356_inw1 = ~( N6809 & N5762 );
	assign N6812 = ~N5762;
	assign AND3_2191_inw1 = ~( N6083 & N6079 );
	assign AND3_2385_inw1 = ~( N6079 & N7191 );
	assign N7188 = ~N6079;
	assign AND3_2384_inw1 = ~( N7188 & N6083 );
	assign N7191 = ~N6083;
	assign N8483 = ~( AND3_2191_inw1 | N6087 );
	assign N8484 = ~( AND3_2192_inw1 | N6087 );
	assign N8469 = ~N6087;
	assign N10062 = ~( N4997 & N9947 );
	assign N6102 = ~N4997;
	assign AND3_2251_inw1 = ~( N6170 & N6166 );
	assign AND3_2395_inw1 = ~( N6166 & N7381 );
	assign N7378 = ~N6166;
	assign AND3_2394_inw1 = ~( N7378 & N6170 );
	assign N7381 = ~N6170;
	assign N8578 = ~( AND3_2251_inw1 | N6174 );
	assign N8579 = ~( AND3_2252_inw1 | N6174 );
	assign N8564 = ~N6174;
	assign N8232 = ~( N6266 & N7580 );
	assign N7581 = ~N6266;
	assign N8233 = ~( N6263 & N7581 );
	assign N7580 = ~N6263;
	assign AND3_2531_inw1 = ~( N6131 & N6127 );
	assign AND3_2636_inw1 = ~( N6127 & N7328 );
	assign N7325 = ~N6127;
	assign N8553 = ~( AND4_2240_inw1 | AND4_2240_inw2 );
	assign AND3_2635_inw1 = ~( N7325 & N6131 );
	assign N7328 = ~N6131;
	assign n_349 = ( N7373 & N7369 );
	assign AND4_2240_inw1 = ~( N7369 & N7358 );
	assign g50_inw1 = ~( N7369 & N7364 );
	assign g58_inw1 = ~( N8552 | N8553 );
	assign N9398 = ~( AND3_2531_inw1 | N7331 );
	assign N9399 = ~( AND3_2532_inw1 | N7331 );
	assign N9394 = ~N7331;
	assign g67_inw1 = ~( N7364 & N7358 );
	assign g55_inw2 = ~( N8418 | n_343 );
	assign AND4_2155_inw1 = ~( N7091 & N7080 );
	assign g48_inw2 = ~( N7080 & n_340 );
	assign g63_inw1 = ~( N7086 & N7080 );
	assign N9396 = ~( AND3_2529_inw1 | N7322 );
	assign N9397 = ~( AND3_2530_inw1 | N7322 );
	assign N9392 = ~N7322;
	assign N8411 = ~( AND4_2151_inw1 | AND4_2151_inw2 );
	assign N8218 = ~( N6246 & N7558 );
	assign N7559 = ~N6246;
	assign AND4_2148_inw1 = ~( N7098 & N7077 );
	assign AND4_2151_inw1 = ~( N7077 & N7068 );
	assign OR4_2378_inw2 = ~( N8410 | N8411 );
	assign N8219 = ~( N6243 & N7559 );
	assign N7558 = ~N6243;
	assign AND4_2148_inw2 = ~( N7073 & N7068 );
	assign g53_inw1 = ~( N7073 & N7068 );
	assign N8950 = ~( OR4_2378_inw1 & OR4_2378_inw2 );
	assign g58_inw2 = ~( N8554 | n_344 );
	assign g50_inw2 = ~( N7358 & n_341 );
	assign N8547 = ~( AND4_2236_inw1 | AND4_2236_inw2 );
	assign AND4_2233_inw1 = ~( N7376 & N7355 );
	assign N9159 = ~( N7577 & N8733 );
	assign N8734 = ~N7577;
	assign AND4_2236_inw1 = ~( N7355 & N7346 );
	assign OR4_2392_inw2 = ~( N8546 | N8547 );
	assign AND4_2233_inw2 = ~( N7351 & N7346 );
	assign g56_inw1 = ~( N7351 & N7346 );
	assign N9160 = ~( N7574 & N8734 );
	assign N8733 = ~N7574;
	assign N9029 = ~( OR4_2392_inw1 & OR4_2392_inw2 );
	assign N9371 = ~( AND3_2517_inw1 | N7213 );
	assign N9372 = ~( AND3_2518_inw1 | N7213 );
	assign N9365 = ~N7213;
	assign N9181 = ~( N7569 & N8755 );
	assign N8756 = ~N7569;
	assign N9182 = ~( N7566 & N8756 );
	assign N8755 = ~N7566;
	assign AND3_2529_inw1 = ~( N7318 & N7314 );
	assign AND3_2634_inw1 = ~( N7314 & N8522 );
	assign N8519 = ~N7314;
	assign n_340 = ( N7099 & N7095 );
	assign N8417 = ~( AND4_2155_inw1 | AND4_2155_inw2 );
	assign n_347 = ( N7095 & N7091 );
	assign AND3_2633_inw1 = ~( N8519 & N7318 );
	assign N8522 = ~N7318;
	assign g48_inw1 = ~( N7091 & N7086 );
	assign g55_inw1 = ~( N8416 | N8417 );
	assign AND3_2515_inw1 = ~( N7198 & N7194 );
	assign AND3_2628_inw1 = ~( N7194 & N8460 );
	assign N8457 = ~N7194;
	assign AND3_2627_inw1 = ~( N8457 & N7198 );
	assign N8460 = ~N7198;
	assign N9369 = ~( AND3_2515_inw1 | N7202 );
	assign N9370 = ~( AND3_2516_inw1 | N7202 );
	assign N9363 = ~N7202;
	assign AND3_2517_inw1 = ~( N7209 & N7205 );
	assign AND3_2630_inw1 = ~( N7205 & N8466 );
	assign N8463 = ~N7205;
	assign AND3_2629_inw1 = ~( N8463 & N7209 );
	assign N8466 = ~N7209;
	assign N9179 = ~( N7563 & N8753 );
	assign N8754 = ~N7563;
	assign N9180 = ~( N7560 & N8754 );
	assign N8753 = ~N7560;
	assign AND3_2547_inw1 = ~( N7398 & N7394 );
	assign AND3_2643_inw1 = ~( N7394 & N8561 );
	assign N8558 = ~N7394;
	assign AND3_2642_inw1 = ~( N8558 & N7398 );
	assign N8561 = ~N7398;
	assign N9421 = ~( AND3_2547_inw1 | N7402 );
	assign N9422 = ~( AND3_2548_inw1 | N7402 );
	assign N9415 = ~N7402;
	assign N9234 = ~( N7591 & N8814 );
	assign N8815 = ~N7591;
	assign N9235 = ~( N7588 & N8815 );
	assign N8814 = ~N7588;
	assign AND3_2545_inw1 = ~( N7387 & N6177 );
	assign AND3_2641_inw1 = ~( N6177 & N8555 );
	assign N7384 = ~N6177;
	assign AND3_2640_inw1 = ~( N7384 & N7387 );
	assign N8555 = ~N7387;
	assign N9419 = ~( AND3_2545_inw1 | N7391 );
	assign N9420 = ~( AND3_2546_inw1 | N7391 );
	assign N9413 = ~N7391;
	assign N9236 = ~( N7585 & N8816 );
	assign N8817 = ~N7585;
	assign N9237 = ~( N7582 & N8817 );
	assign N8816 = ~N7582;
	assign N9146 = ~NOR3_2424_invw;
	assign N10195 = ~N9979;
	assign N10892 = ~( N10857 & N10816 );
	assign N10950 = ~( N10919 & N10891 );
	assign N10816 = ~( N10691 & N9741 );
	assign N10891 = ~( N10812 & N9741 );
	assign N10333 = ~( N10192 & N9977 );
	assign N10332 = ~N10192;
	assign N10759 = ( N10705 | N10549 );
	assign N10706 = ( N10631 | N10551 );
	assign N9837 = ~N9429;
	assign N6191 = ~N4784;
	assign g3_inw2 = ~( n_316 | n_317 );
	assign g73_inw2 = ~( n_316 | n_352 );
	assign N9426 = ~( N9064 & N8608 );
	assign N10837 = ( N10730 | N10587 );
	assign N10546 = ( N5631 & N10450 );
	assign N10102 = ~( g32_inw1 & g32_inw2 );
	assign N9736 = ( N9265 & N8262 );
	assign N10020 = ~( AND3_2834_inw1 | N8262 );
	assign AND4_2835_inw2 = ~( N8298 & N8262 );
	assign N9732 = ( N9265 & N8269 );
	assign N10013 = ~( AND3_2827_inw1 | N8269 );
	assign AND4_2828_inw2 = ~( N8307 & N8269 );
	assign AND3_3101_inw1 = ~( N10357 & N9905 );
	assign AND3_3132_inw1 = ~( N10357 & N7609 );
	assign AND3_3100_inw1 = ~( N10360 & N9543 );
	assign AND3_3131_inw1 = ~( N10360 & N8857 );
	assign N10840 = N10839;
	assign N10241 = ~N10070;
	assign N10242 = ~N10073;
	assign N9526 = ( N8943 & N8421 );
	assign N10016 = ~( AND3_2830_inw1 | N8421 );
	assign AND4_2831_inw2 = ~( N8394 & N8421 );
	assign N10587 = ( N10367 & N5735 );
	assign N10234 = ~( N7100 & N10140 );
	assign N10295 = ~( N8412 & N10233 );
	assign N11213 = ~N11168;
	assign N11215 = ~N11171;
	assign N10282 = ( N6784 & N10141 );
	assign N10270 = ~( N6762 & N10116 );
	assign N8254 = ~N6762;
	assign N7609 = ~( g7_inw1 & g7_inw2 );
	assign N8131 = ~NOR3_2032_invw;
	assign N9066 = ~N8114;
	assign N10568 = ~N10422;
	assign N10647 = ~( AND3_3130_inw1 | N10577 );
	assign N10076 = ~( N9068 & N9957 );
	assign N9645 = ~N9068;
	assign N10872 = ~N10789;
	assign N10874 = ~N10792;
	assign N9959 = ~N9646;
	assign N9958 = ~( N9642 & N9645 );
	assign N9957 = ~N9642;
	assign N10570 = ~N10425;
	assign N10988 = ~N10928;
	assign N10990 = ~N10931;
	assign N10173 = ~( N10077 & N9960 );
	assign N10077 = ~( N9074 & N9959 );
	assign N10419 = ~( g93_inw1 & g93_inw2 );
	assign N8117 = ~( g103_inw1 & g103_inw2 );
	assign N11278 = ( N10116 & N11260 );
	assign N11277 = ~N11261;
	assign N8134 = ~NOR4_2033_invw;
	assign N11114 = ~N11044;
	assign N11116 = ~N11047;
	assign N10082 = ~( N9089 & N9967 );
	assign N9666 = ~N9089;
	assign N10882 = ~N10800;
	assign N10884 = ~N10803;
	assign N8183 = ~NOR3_2040_invw;
	assign N9969 = ~N9667;
	assign N9968 = ~( N9663 & N9666 );
	assign N9967 = ~N9663;
	assign N10561 = ~N10412;
	assign N10998 = ~N10938;
	assign N11000 = ~N10941;
	assign N8307 = ( N6833 & N6881 );
	assign N10183 = ~( N10083 & N9970 );
	assign N10083 = ~( N9095 & N9969 );
	assign N11217 = ~N11174;
	assign N11219 = ~N11177;
	assign N8298 = ( N6833 & N6845 );
	assign N8288 = ~N6845;
	assign N7655 = ~( g19_inw1 & g19_inw2 );
	assign N9087 = ~N8166;
	assign N10559 = ~N10409;
	assign N10406 = ~( g89_inw1 & g89_inw2 );
	assign N8169 = ~( g101_inw1 & g101_inw2 );
	assign N11279 = ~N11263;
	assign N8186 = ~NOR4_2041_invw;
	assign N11118 = ~N11050;
	assign N11120 = ~N11053;
	assign N9659 = ~N9079;
	assign N8883 = ~N8204;
	assign N8874 = ( N6833 & N7655 );
	assign N10796 = ~N10675;
	assign N10798 = ~N10678;
	assign N10709 = ( N9243 & N10589 );
	assign N10179 = ~( N9964 & N8881 );
	assign N10178 = ~N9964;
	assign N9541 = ~N9275;
	assign N10177 = ~( N9961 & N8879 );
	assign N10176 = ~N9961;
	assign N10934 = ~N10876;
	assign N10936 = ~N10879;
	assign N8156 = ~NOR3_2037_invw;
	assign N10554 = ( N10375 & N9540 );
	assign N9738 = ~N9556;
	assign AND3_3403_inw1 = ~( N11100 & N7655 );
	assign AND3_3405_inw1 = ~( N11100 & N9917 );
	assign AND3_3402_inw1 = ~( N11103 & N8871 );
	assign AND3_3404_inw1 = ~( N11103 & N9551 );
	assign N10247 = ~( N8146 & N10176 );
	assign N8879 = ~N8146;
	assign N10553 = ( N10375 & N9539 );
	assign N9737 = ~N9555;
	assign N11040 = ~N10992;
	assign N11042 = ~N10995;
	assign N9265 = ( N7649 | N8874 );
	assign N10441 = ~( N9682 & N10332 );
	assign N9977 = ~N9682;
	assign N11065 = ~N11008;
	assign N11122 = ~N11062;
	assign N9754 = ( N8333 & N9280 );
	assign N10334 = ~( N10259 & N10196 );
	assign N10259 = ~( N9692 & N10195 );
	assign N11264 = ~N11233;
	assign N11290 = ~N11272;
	assign N9775 = ( N8333 & N9307 );
	assign N9769 = ~N9307;
	assign N8902 = ~( g23_inw1 & g23_inw2 );
	assign N9899 = ~N9629;
	assign N9975 = ~N9679;
	assign N9626 = ~( g85_inw1 & g85_inw2 );
	assign N9685 = ~( g107_inw1 & g107_inw2 );
	assign N11296 = ~N11292;
	assign N9149 = ~NOR4_2425_invw;
	assign N11183 = ~N11124;
	assign N11231 = ~N11180;
	assign N9971 = ~N9671;
	assign N9565 = ~N9107;
	assign N9560 = ( N8902 & N8333 );
	assign N9276 = ~N8333;
	assign N10886 = ~N10806;
	assign N10888 = ~N10809;
	assign N10331 = ~( N10189 & N9563 );
	assign N10330 = ~N10189;
	assign N9896 = ~N9766;
	assign N10329 = ~( N10186 & N9561 );
	assign N10328 = ~N10186;
	assign N11002 = ~N10944;
	assign N11004 = ~N10947;
	assign N9103 = ~NOR3_2419_invw;
	assign N10028 = ~N9924;
	assign AND3_3434_inw1 = ~( N11156 & N8902 );
	assign AND3_3436_inw1 = ~( N11156 & N10132 );
	assign AND3_3433_inw1 = ~( N11159 & N9575 );
	assign AND3_3435_inw1 = ~( N11159 & N9935 );
	assign N10439 = ~( N9099 & N10328 );
	assign N9561 = ~N9099;
	assign N10026 = ~N9923;
	assign N11106 = ~N11056;
	assign N11108 = ~N11059;
	assign N9557 = ~N8898;
	assign N9758 = ( N8898 | N9560 );
	assign N10264 = ~( N9717 & N10203 );
	assign N10002 = ~N9717;
	assign N10961 = ~N10899;
	assign N10963 = ~N10902;
	assign N9220 = ~NOR3_2440_invw;
	assign N10205 = ~N10003;
	assign N10204 = ~( N9999 & N10002 );
	assign N10203 = ~N9999;
	assign N10773 = ~N10665;
	assign N11073 = ~N11015;
	assign N11075 = ~N11018;
	assign N9344 = ( N8430 & N8444 );
	assign N10598 = ( N8444 & N10381 );
	assign N10344 = ~( N10265 & N10206 );
	assign N10265 = ~( N9723 & N10205 );
	assign N11267 = ~N11236;
	assign N11269 = ~N11239;
	assign N9385 = ( N8430 & N8497 );
	assign N9375 = ~N8497;
	assign N8966 = ~( g21_inw1 & g21_inw2 );
	assign N9715 = ~N9203;
	assign N10771 = ~N10662;
	assign N10659 = ~( g97_inw1 & g97_inw2 );
	assign N9206 = ~( g105_inw1 & g105_inw2 );
	assign N11298 = ( N10301 & N11293 );
	assign N11297 = ~N11294;
	assign N9223 = ~NOR4_2441_invw;
	assign N11185 = ~N11127;
	assign N11187 = ~N11130;
	assign N9995 = ~N9707;
	assign N9596 = ~N9169;
	assign N9591 = ( N8966 & N8430 );
	assign N10895 = ~N10817;
	assign N10897 = ~N10820;
	assign N10866 = ( N9739 & N10784 );
	assign N10340 = ~( N10200 & N9594 );
	assign N10339 = ~N10200;
	assign N9892 = ~N9799;
	assign N10338 = ~( N10197 & N9592 );
	assign N10337 = ~N10197;
	assign N11011 = ~N10955;
	assign N11013 = ~N10958;
	assign N9165 = ~NOR3_2429_invw;
	assign N10766 = ( N10652 & N9891 );
	assign N10024 = ~N9946;
	assign AND3_3438_inw1 = ~( N11162 & N8966 );
	assign AND3_3440_inw1 = ~( N11162 & N10160 );
	assign AND3_3437_inw1 = ~( N11165 & N9608 );
	assign AND3_3439_inw1 = ~( N11165 & N9949 );
	assign N10444 = ~( N9161 & N10337 );
	assign N9592 = ~N9161;
	assign N10765 = ( N10652 & N9890 );
	assign N10023 = ~N9945;
	assign N11110 = ~N11067;
	assign N11112 = ~N11070;
	assign N9791 = ( N8963 | N9591 );
	assign N10719 = ~N10381;
	assign N11342 = ~N11341;
	assign N11302 = ( N11289 | N11280 );
	assign OR4_3421_inw2 = ~( N11154 | N11155 );
	assign N11289 = ( N11279 & N10283 );
	assign N11152 = ~( AND3_3402_inw1 | N10283 );
	assign N11153 = ~( AND3_3403_inw1 | N10283 );
	assign N10375 = ( N7655 | N10291 );
	assign N10581 = ~( AND3_3100_inw1 | N10116 );
	assign N10582 = ~( AND3_3101_inw1 | N10116 );
	assign N10479 = ~N10116;
	assign N10465 = ~N10141;
	assign N11228 = ~( AND3_3439_inw1 | N10301 );
	assign N11229 = ~( AND3_3440_inw1 | N10301 );
	assign N10497 = ~N10301;
	assign N10101 = ~( g3_inw1 & g3_inw2 );
	assign N10104 = ~( g73_inw1 & g73_inw2 );
	assign N8863 = ~( AND3_2354_inw1 | N8276 );
	assign N7100 = ~( g46_inw1 | g46_inw2 );
	assign N9258 = ~( N8863 | N8282 );
	assign N9259 = ~( N8864 | N8283 );
	assign N7826 = ~( g52_inw1 & g52_inw2 );
	assign N8394 = ~( g39_inw1 | g39_inw2 );
	assign N9400 = ~( N9024 | N8539 );
	assign N9401 = ~( N9025 | N8540 );
	assign N9024 = ~( AND3_2390_inw1 | N8537 );
	assign N9025 = ~( AND3_2391_inw1 | N8537 );
	assign N7057 = ~( AND4_1866_inw1 | AND4_1866_inw2 );
	assign N8727 = ~( N8216 & N8217 );
	assign N8943 = ( N7825 | N8404 );
	assign N9260 = ~( N8865 | N8284 );
	assign N9261 = ~( N8866 | N8285 );
	assign N8865 = ~( AND3_2356_inw1 | N8278 );
	assign N8866 = ~( AND3_2357_inw1 | N8278 );
	assign N8627 = ~( N8144 & N8145 );
	assign N8861 = ~( AND3_2352_inw1 | N8274 );
	assign N9256 = ~( N8861 | N8280 );
	assign N9257 = ~( N8862 | N8281 );
	assign N10113 = ~( N10036 & N9907 );
	assign N9907 = ~( N9650 & N5769 );
	assign N10114 = ~( N10037 & N9909 );
	assign N9909 = ~( N9653 & N5770 );
	assign N8959 = ~N7852;
	assign AND3_2232_inw1 = ~( N7337 & N7334 );
	assign g39_inw2 = ~( n_335 & n_336 );
	assign AND3_2080_inw1 = ~( N6812 & N6809 );
	assign N8992 = ~( AND3_2385_inw1 | N8469 );
	assign AND3_2192_inw1 = ~( N7191 & N7188 );
	assign N8991 = ~( AND3_2384_inw1 | N8469 );
	assign N9367 = ~( N8991 | N8483 );
	assign N9368 = ~( N8992 | N8484 );
	assign N10155 = ~( N10062 & N9948 );
	assign N9948 = ~( N9702 & N6102 );
	assign N9054 = ~( AND3_2395_inw1 | N8564 );
	assign AND3_2252_inw1 = ~( N7381 & N7378 );
	assign N9053 = ~( AND3_2394_inw1 | N8564 );
	assign N9417 = ~( N9053 | N8578 );
	assign N9418 = ~( N9054 | N8579 );
	assign N8811 = ~( N8232 & N8233 );
	assign N9615 = ~( AND3_2636_inw1 | N9394 );
	assign AND3_2532_inw1 = ~( N7328 & N7325 );
	assign N9614 = ~( AND3_2635_inw1 | N9394 );
	assign N8548 = ~( g50_inw1 | g50_inw2 );
	assign N9035 = ~( g58_inw1 & g58_inw2 );
	assign N9815 = ~( N9614 | N9398 );
	assign N9816 = ~( N9615 | N9399 );
	assign N8956 = ~( g55_inw1 & g55_inw2 );
	assign N8412 = ~( g48_inw1 | g48_inw2 );
	assign N9813 = ~( N9612 | N9396 );
	assign N9814 = ~( N9613 | N9397 );
	assign N9612 = ~( AND3_2633_inw1 | N9392 );
	assign N9613 = ~( AND3_2634_inw1 | N9392 );
	assign N8730 = ~( N8218 & N8219 );
	assign N8405 = ~( AND4_2148_inw1 | AND4_2148_inw2 );
	assign N10548 = ( N10391 & N8950 );
	assign N9581 = ~N8950;
	assign N9786 = ( N8950 | N9585 );
	assign N8541 = ~( AND4_2233_inw1 | AND4_2233_inw2 );
	assign N9478 = ~( N9159 & N9160 );
	assign N9616 = ~N9029;
	assign N9820 = ( N9029 | N9618 );
	assign N9802 = ~( N9604 | N9371 );
	assign N9803 = ~( N9605 | N9372 );
	assign N9604 = ~( AND3_2629_inw1 | N9365 );
	assign N9605 = ~( AND3_2630_inw1 | N9365 );
	assign N9488 = ~( N9181 & N9182 );
	assign AND3_2530_inw1 = ~( N8522 & N8519 );
	assign N9603 = ~( AND3_2628_inw1 | N9363 );
	assign AND3_2516_inw1 = ~( N8460 & N8457 );
	assign N9602 = ~( AND3_2627_inw1 | N9363 );
	assign N9800 = ~( N9602 | N9369 );
	assign N9801 = ~( N9603 | N9370 );
	assign AND3_2518_inw1 = ~( N8466 & N8463 );
	assign N9485 = ~( N9179 & N9180 );
	assign N9624 = ~( AND3_2643_inw1 | N9415 );
	assign AND3_2548_inw1 = ~( N8561 & N8558 );
	assign N9623 = ~( AND3_2642_inw1 | N9415 );
	assign N9829 = ~( N9623 | N9421 );
	assign N9830 = ~( N9624 | N9422 );
	assign N9517 = ~( N9234 & N9235 );
	assign N9622 = ~( AND3_2641_inw1 | N9413 );
	assign AND3_2546_inw1 = ~( N8555 & N7384 );
	assign N9621 = ~( AND3_2640_inw1 | N9413 );
	assign N9827 = ~( N9621 | N9419 );
	assign N9828 = ~( N9622 | N9420 );
	assign N9520 = ~( N9236 & N9237 );
	assign N9690 = ~N9146;
	assign N10953 = ~N10892;
	assign N11006 = ~N10950;
	assign N10531 = ~( N10441 & N10333 );
	assign N9835 = ~N9426;
	assign N10838 = N10837;
	assign N10103 = N10102;
	assign n_352 = ( N9736 | N10020 );
	assign N10021 = ~( AND4_2835_inw1 | AND4_2835_inw2 );
	assign n_317 = ( N9732 | N10013 );
	assign N10014 = ~( AND4_2828_inw1 | AND4_2828_inw2 );
	assign N10649 = ~( AND3_3132_inw1 | N10479 );
	assign N10648 = ~( AND3_3131_inw1 | N10479 );
	assign n_332 = ( N9526 | N10016 );
	assign N10017 = ~( AND4_2831_inw1 | AND4_2831_inw2 );
	assign N10296 = ( N8959 & N10234 );
	assign N10391 = ( N9582 & N10295 );
	assign N10367 = ( N7609 | N10282 );
	assign N10354 = ( N8857 & N10270 );
	assign N9543 = ( N8857 & N8254 );
	assign N8857 = ~N7609;
	assign N9072 = ~N8131;
	assign N10729 = ~N10647;
	assign N10170 = ~( N10076 & N9958 );
	assign N10317 = ~( N10173 & N9077 );
	assign N10316 = ~N10173;
	assign N10566 = ~N10419;
	assign N10431 = ~( N8117 & N10314 );
	assign N9071 = ~N8117;
	assign N11299 = ( N11288 | N11278 );
	assign N11288 = ( N11277 & N10479 );
	assign N10432 = ~( N8134 & N10316 );
	assign N9077 = ~N8134;
	assign N10180 = ~( N10082 & N9968 );
	assign N9093 = ~N8183;
	assign N10057 = ( N9791 & N8307 );
	assign AND3_2827_inw1 = ~( N9791 & N8307 );
	assign N10058 = ~( AND3_2860_inw1 | N8307 );
	assign AND4_2861_inw2 = ~( N9344 & N8307 );
	assign g5_inw1 = ~( N9344 & N8307 );
	assign N10327 = ~( N10183 & N9098 );
	assign N10326 = ~N10183;
	assign N10039 = ( N9791 & N8298 );
	assign AND3_2834_inw1 = ~( N9791 & N8298 );
	assign N10040 = ~( AND3_2850_inw1 | N8298 );
	assign AND4_2851_inw2 = ~( N9385 & N8298 );
	assign g75_inw1 = ~( N9385 & N8298 );
	assign N9551 = ( N8871 & N8288 );
	assign N8871 = ~N7655;
	assign N10557 = ~N10406;
	assign N10437 = ~( N8169 & N10324 );
	assign N9092 = ~N8169;
	assign N10438 = ~( N8186 & N10326 );
	assign N9098 = ~N8186;
	assign N10762 = ( N10709 | N10555 );
	assign N10321 = ~( N10248 & N10179 );
	assign N10248 = ~( N8156 & N10178 );
	assign N10555 = ( N10375 & N9541 );
	assign N10318 = ~( N10247 & N10177 );
	assign N8881 = ~N8156;
	assign N10761 = ( N10708 | N10554 );
	assign N10708 = ( N9738 & N10589 );
	assign N10760 = ( N10707 | N10553 );
	assign N10707 = ( N9737 & N10589 );
	assign OR4_2892_inw1 = ~( N9265 | N10039 );
	assign OR4_2906_inw1 = ~( N9265 | N10057 );
	assign N10535 = ~( N10334 & N9695 );
	assign N10534 = ~N10334;
	assign N9935 = ( N9575 & N9769 );
	assign N9575 = ~N8902;
	assign N9897 = ~N9626;
	assign N10750 = ~( N9685 & N10689 );
	assign N9978 = ~N9685;
	assign N10621 = ~( N9149 & N10534 );
	assign N9695 = ~N9149;
	assign N9768 = ~( N9557 & N9276 );
	assign N10528 = ~( N10440 & N10331 );
	assign N10440 = ~( N9103 & N10330 );
	assign N10525 = ~( N10439 & N10329 );
	assign N9563 = ~N9103;
	assign N10042 = ( N9758 & N9385 );
	assign N10060 = ( N9758 & N9344 );
	assign AND3_2850_inw1 = ~( N9758 & N9385 );
	assign AND3_2860_inw1 = ~( N9758 & N9344 );
	assign AND4_2828_inw1 = ~( N9758 & N9344 );
	assign AND4_2835_inw1 = ~( N9758 & N9385 );
	assign N10341 = ~( N10264 & N10204 );
	assign N9721 = ~N9220;
	assign N10652 = ( N8966 | N10598 );
	assign N10545 = ~( N10344 & N9726 );
	assign N10544 = ~N10344;
	assign N9949 = ( N9608 & N9375 );
	assign N9608 = ~N8966;
	assign N10769 = ~N10659;
	assign N10626 = ~( N9206 & N10542 );
	assign N9720 = ~N9206;
	assign N11317 = ( N11309 | N11298 );
	assign N11309 = ( N11297 & N10497 );
	assign N10627 = ~( N9223 & N10544 );
	assign N9726 = ~N9223;
	assign N10907 = ( N10866 | N10767 );
	assign N10539 = ~( N10445 & N10340 );
	assign N10445 = ~( N9165 & N10339 );
	assign N10767 = ( N10652 & N9892 );
	assign N10536 = ~( N10444 & N10338 );
	assign N9594 = ~N9165;
	assign N10906 = ( N10865 | N10766 );
	assign N10865 = ( N10024 & N10784 );
	assign N11227 = ~( AND3_3438_inw1 | N10497 );
	assign N11226 = ~( AND3_3437_inw1 | N10497 );
	assign N10905 = ( N10864 | N10765 );
	assign N10864 = ( N10023 & N10784 );
	assign OR3_2893_inw1 = ~( N9791 | N10042 );
	assign OR3_2907_inw1 = ~( N9791 | N10060 );
	assign N11312 = ~( N11302 & N11246 );
	assign N11315 = ~N11302;
	assign N11205 = ~( OR4_3421_inw1 & OR4_3421_inw2 );
	assign OR4_3421_inw1 = ~( N11152 | N11153 );
	assign N10589 = ~N10375;
	assign OR4_3183_inw2 = ~( N10581 | N10582 );
	assign OR4_3453_inw2 = ~( N11228 | N11229 );
	assign N9653 = ~( N9259 & N9258 );
	assign N8404 = ( N7057 & N7826 );
	assign N10055 = ( N9786 & N8394 );
	assign AND3_2830_inw1 = ~( N9786 & N8394 );
	assign N10056 = ~( AND3_2858_inw1 | N8394 );
	assign AND4_2717_inw2 = ~( N9332 & N8394 );
	assign g34_inw1 = ~( N9332 & N8394 );
	assign N9698 = ~( N9401 & N9400 );
	assign N10050 = ~( N8727 & N9938 );
	assign N9323 = ~N8727;
	assign OR4_2905_inw1 = ~( N8943 | N10055 );
	assign N9656 = ~( N9261 & N9260 );
	assign N10038 = ~( N8627 & N9910 );
	assign N9262 = ~N8627;
	assign N9650 = ~( N9257 & N9256 );
	assign AND4_3022_inw1 = ~( N10113 & N10115 );
	assign AND4_3020_inw1 = ~( N10114 & N10134 );
	assign N9702 = ~( N9368 & N9367 );
	assign AND4_3023_inw1 = ~( N10155 & N10161 );
	assign N9727 = ~( N9418 & N9417 );
	assign N10067 = ~( N8811 & N9953 );
	assign N9412 = ~N8811;
	assign N9408 = ( N8541 & N8548 );
	assign N9618 = ( N8541 & N9035 );
	assign N9617 = ~N9035;
	assign N9986 = ~( N9816 & N9815 );
	assign N9585 = ( N8405 & N8956 );
	assign N9582 = ~N8956;
	assign N9332 = ( N8405 & N8412 );
	assign N9983 = ~( N9814 & N9813 );
	assign N10231 = ~( N8730 & N10135 );
	assign N9324 = ~N8730;
	assign N9326 = ~N8405;
	assign N10704 = ( N10629 | N10548 );
	assign N9733 = ~( N9581 & N9326 );
	assign N9402 = ~N8541;
	assign N10232 = ~( N9478 & N10137 );
	assign N9784 = ~N9478;
	assign N9785 = ~( N9616 & N9402 );
	assign AND3_2858_inw1 = ~( N9820 & N9332 );
	assign AND4_2831_inw1 = ~( N9820 & N9332 );
	assign N9992 = ~( N9803 & N9802 );
	assign N10238 = ~( N9488 & N10158 );
	assign N9806 = ~N9488;
	assign N9989 = ~( N9801 & N9800 );
	assign N10237 = ~( N9485 & N10156 );
	assign N9805 = ~N9485;
	assign N10007 = ~( N9830 & N9829 );
	assign N10239 = ~( N9517 & N10162 );
	assign N9825 = ~N9517;
	assign N10010 = ~( N9828 & N9827 );
	assign N10240 = ~( N9520 & N10164 );
	assign N9826 = ~N9520;
	assign N10690 = ~( N10531 & N9978 );
	assign N10689 = ~N10531;
	assign OR4_3183_inw1 = ~( N10648 | N10649 );
	assign N10450 = ~N10296;
	assign N10547 = ~N10391;
	assign N10583 = ~N10367;
	assign N10550 = ~N10354;
	assign N9905 = ~N9543;
	assign N10315 = ~( N10170 & N9071 );
	assign N10314 = ~N10170;
	assign N10512 = ~( N10432 & N10317 );
	assign N10509 = ~( N10431 & N10315 );
	assign N11313 = ~( N11299 & N10836 );
	assign N11314 = ~N11299;
	assign N10325 = ~( N10180 & N9092 );
	assign N10324 = ~N10180;
	assign N10522 = ~( N10438 & N10327 );
	assign N9917 = ~N9551;
	assign N10519 = ~( N10437 & N10325 );
	assign N10517 = ~N10321;
	assign N10515 = ~N10318;
	assign N10691 = ~( N10621 & N10535 );
	assign N10132 = ~N9935;
	assign N10812 = ~( N10750 & N10690 );
	assign N10687 = ~N10528;
	assign N10685 = ~N10525;
	assign N10543 = ~( N10341 & N9720 );
	assign N10542 = ~N10341;
	assign N10784 = ~N10652;
	assign N10701 = ~( N10627 & N10545 );
	assign N10160 = ~N9949;
	assign N10698 = ~( N10626 & N10543 );
	assign N11329 = ~( N11317 & N11286 );
	assign N11331 = ~N11317;
	assign N10696 = ~N10539;
	assign N10694 = ~N10536;
	assign OR4_3453_inw1 = ~( N11226 | N11227 );
	assign N11327 = ~( N11312 & N11320 );
	assign N11320 = ~( N11205 & N11315 );
	assign N11246 = ~N11205;
	assign N10739 = ~( OR4_3183_inw1 & OR4_3183_inw2 );
	assign N11257 = ~( OR4_3453_inw1 & OR4_3453_inw2 );
	assign N9908 = ~N9653;
	assign N9939 = ~( N9698 & N9323 );
	assign N9938 = ~N9698;
	assign N10134 = ~( N10050 & N9939 );
	assign N9911 = ~( N9656 & N9262 );
	assign N9910 = ~N9656;
	assign N10115 = ~( N10038 & N9911 );
	assign N9906 = ~N9650;
	assign N10399 = ~( AND4_3022_inw1 | AND4_3022_inw2 );
	assign N10388 = ~( AND4_3020_inw1 | AND4_3020_inw2 );
	assign N9947 = ~N9702;
	assign N10402 = ~( AND4_3023_inw1 | AND4_3023_inw2 );
	assign N9954 = ~( N9727 & N9412 );
	assign N9953 = ~N9727;
	assign N10161 = ~( N10067 & N9954 );
	assign N10138 = ~( N9986 & N9784 );
	assign N10137 = ~N9986;
	assign N10136 = ~( N9983 & N9324 );
	assign N10135 = ~N9983;
	assign N10293 = ~( N10231 & N10136 );
	assign N10629 = ( N9733 & N10547 );
	assign N10294 = ~( N10232 & N10138 );
	assign N10159 = ~( N9992 & N9806 );
	assign N10158 = ~N9992;
	assign N10300 = ~( N10238 & N10159 );
	assign N10157 = ~( N9989 & N9805 );
	assign N10156 = ~N9989;
	assign N10299 = ~( N10237 & N10157 );
	assign N10163 = ~( N10007 & N9825 );
	assign N10162 = ~N10007;
	assign N10306 = ~( N10239 & N10163 );
	assign N10165 = ~( N10010 & N9826 );
	assign N10164 = ~N10010;
	assign N10307 = ~( N10240 & N10165 );
	assign N10673 = ~N10512;
	assign N10671 = ~N10509;
	assign N11328 = ~( N11313 & N11321 );
	assign N11321 = ~( N10739 & N11314 );
	assign N10683 = ~N10522;
	assign N10681 = ~N10519;
	assign N10815 = ~N10691;
	assign N10890 = ~N10812;
	assign N10825 = ~N10701;
	assign N10823 = ~N10698;
	assign N11338 = ~( N11329 & N11335 );
	assign N11335 = ~( N11257 & N11331 );
	assign N11333 = ~N11327;
	assign N10836 = ~N10739;
	assign N11286 = ~N11257;
	assign AND3_3099_inw1 = ~( N10399 & N10402 );
	assign N10574 = ~N10399;
	assign N10577 = ~( AND3_3099_inw1 | N10388 );
	assign N10576 = ~N10388;
	assign N10575 = ~N10402;
	assign AND4_3020_inw2 = ~( N10293 & N10294 );
	assign AND4_3022_inw2 = ~( N10299 & N10300 );
	assign AND4_3023_inw2 = ~( N10306 & N10307 );
	assign N11334 = ~N11328;
	assign N11340 = ~N11338;
endmodule
